// soc_system.v

// Generated using ACDS version 13.1 162 at 2014.12.19.15:54:10

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                                  //                         clk.clk
		input  wire        reset_reset_n,                            //                       reset.reset_n
		output wire [14:0] memory_mem_a,                             //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                            //                            .mem_ba
		output wire        memory_mem_ck,                            //                            .mem_ck
		output wire        memory_mem_ck_n,                          //                            .mem_ck_n
		output wire        memory_mem_cke,                           //                            .mem_cke
		output wire        memory_mem_cs_n,                          //                            .mem_cs_n
		output wire        memory_mem_ras_n,                         //                            .mem_ras_n
		output wire        memory_mem_cas_n,                         //                            .mem_cas_n
		output wire        memory_mem_we_n,                          //                            .mem_we_n
		output wire        memory_mem_reset_n,                       //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                            //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                           //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                         //                            .mem_dqs_n
		output wire        memory_mem_odt,                           //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                            //                            .mem_dm
		input  wire        memory_oct_rzqin,                         //                            .oct_rzqin
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,    //                hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,      //                            .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,      //                            .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,      //                            .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,      //                            .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,      //                            .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,      //                            .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,       //                            .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,    //                            .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,    //                            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,    //                            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,      //                            .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,      //                            .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,      //                            .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,        //                            .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,        //                            .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,        //                            .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,        //                            .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,        //                            .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,        //                            .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,        //                            .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,         //                            .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,         //                            .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,        //                            .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,         //                            .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,         //                            .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,         //                            .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,         //                            .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,         //                            .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,         //                            .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,         //                            .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,         //                            .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,         //                            .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,         //                            .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,        //                            .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,        //                            .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,        //                            .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,        //                            .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,       //                            .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,      //                            .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,      //                            .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,       //                            .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,        //                            .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,        //                            .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,        //                            .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,        //                            .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,        //                            .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,        //                            .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,     //                            .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,     //                            .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,     //                            .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,     //                            .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,     //                            .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,     //                            .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,     //                            .hps_io_gpio_inst_GPIO61
		output wire        hps_0_h2f_reset_reset_n,                  //             hps_0_h2f_reset.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,     //     hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,         //    hps_0_f2h_warm_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,        //   hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_cold_reset_req_reset_n,         //    hps_0_f2h_cold_reset_req.reset_n
		output wire [1:0]  pio_alivetest_cpu_s0_extcon_export,       // pio_alivetest_cpu_s0_extcon.export
		output wire [12:0] sdram_wire_addr,                          //                  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                            //                            .ba
		output wire        sdram_wire_cas_n,                         //                            .cas_n
		output wire        sdram_wire_cke,                           //                            .cke
		output wire        sdram_wire_cs_n,                          //                            .cs_n
		inout  wire [15:0] sdram_wire_dq,                            //                            .dq
		output wire [1:0]  sdram_wire_dqm,                           //                            .dqm
		output wire        sdram_wire_ras_n,                         //                            .ras_n
		output wire        sdram_wire_we_n,                          //                            .we_n
		output wire [1:0]  pio_alivetest_cpu_s1_extcon_export,       // pio_alivetest_cpu_s1_extcon.export
		output wire        system_pll_locked_export,                 //           system_pll_locked.export
		output wire        sdram_pll_locked_export,                  //            sdram_pll_locked.export
		inout  wire        i2c_cpu_s0_i2c_exports_scl,               //      i2c_cpu_s0_i2c_exports.scl
		inout  wire        i2c_cpu_s0_i2c_exports_sda,               //                            .sda
		inout  wire        i2c_cpu_s1_i2c_exports_scl,               //      i2c_cpu_s1_i2c_exports.scl
		inout  wire        i2c_cpu_s1_i2c_exports_sda,               //                            .sda
		output wire        pwm_cpu_s0_1_conduit_end_readdatavalid_n, //    pwm_cpu_s0_1_conduit_end.readdatavalid_n
		output wire        clk_sdram_clk,                            //                   clk_sdram.clk
		output wire        pwm_cpu_s0_2_conduit_end_readdatavalid_n, //    pwm_cpu_s0_2_conduit_end.readdatavalid_n
		output wire        pwm_cpu_s0_3_conduit_end_readdatavalid_n, //    pwm_cpu_s0_3_conduit_end.readdatavalid_n
		output wire        pwm_cpu_s0_4_conduit_end_readdatavalid_n, //    pwm_cpu_s0_4_conduit_end.readdatavalid_n
		output wire        pwm_cpu_s0_5_conduit_end_readdatavalid_n, //    pwm_cpu_s0_5_conduit_end.readdatavalid_n
		output wire        pwm_cpu_s0_6_conduit_end_readdatavalid_n, //    pwm_cpu_s0_6_conduit_end.readdatavalid_n
		output wire        pwm_cpu_s0_7_conduit_end_readdatavalid_n, //    pwm_cpu_s0_7_conduit_end.readdatavalid_n
		output wire        pwm_cpu_s0_8_conduit_end_readdatavalid_n  //    pwm_cpu_s0_8_conduit_end.readdatavalid_n
	);

	wire         system_pll_outclk0_clk;                                           // system_pll:outclk_0 -> [cpu_s0:clk, cpu_s1:clk, fifo_bridge_cpuM_cpus0:clk, fifo_bridge_cpuM_cpus1:clk, fifo_bridge_cpus0_cpus1:clk, fpga_only_master:clk_clk, hps_only_master:clk_clk, intr_capturer_0:clk, irq_mapper_002:clk, irq_mapper_003:clk, irq_mapper_004:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, irq_synchronizer_005:sender_clk, mm_interconnect_0:system_pll_outclk0_clk, mm_interconnect_1:system_pll_outclk0_clk, mm_interconnect_2:system_pll_outclk0_clk, mm_interconnect_3:system_pll_outclk0_clk, mm_interconnect_4:system_pll_outclk0_clk, onchip_sram:clk, rst_controller:clk, s0_io_clockCrossing_bridge:s0_clk, s1_io_clockCrossing_bridge:s0_clk, sdram_clockCrossing_Bridge:s0_clk, sysid_qsys:clock]
	wire         system_pll_outclk1_clk;                                           // system_pll:outclk_1 -> [i2c_cpu_s0:wb_clk_i, i2c_cpu_s1:wb_clk_i, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, irq_synchronizer_004:receiver_clk, irq_synchronizer_005:receiver_clk, jtag_uart_cpu_s0:clk, jtag_uart_cpu_s1:clk, mm_interconnect_5:system_pll_outclk1_clk, mm_interconnect_7:system_pll_outclk1_clk, pio_aliveTest_cpu_s0:clk, pio_aliveTest_cpu_s1:clk, rst_controller_001:clk, s0_io_clockCrossing_bridge:m0_clk, s1_io_clockCrossing_bridge:m0_clk, timer_cpu_s0:clk, timer_cpu_s1:clk]
	wire         sdram_pll_outclk0_clk;                                            // sdram_pll:outclk_0 -> [mm_interconnect_6:sdram_pll_outclk0_clk, rst_controller_002:clk, sdram:clk, sdram_clockCrossing_Bridge:m0_clk]
	wire         pwm_pll_outclk0_clk;                                              // pwm_pll:outclk_0 -> [mm_interconnect_5:pwm_pll_outclk0_clk, pwm_cpu_s0_1:clk, pwm_cpu_s0_2:clk, pwm_cpu_s0_3:clk, pwm_cpu_s0_4:clk, pwm_cpu_s0_5:clk, pwm_cpu_s0_6:clk, pwm_cpu_s0_7:clk, pwm_cpu_s0_8:clk, rst_controller_004:clk]
	wire         hps_only_master_master_waitrequest;                               // mm_interconnect_0:hps_only_master_master_waitrequest -> hps_only_master:master_waitrequest
	wire  [31:0] hps_only_master_master_writedata;                                 // hps_only_master:master_writedata -> mm_interconnect_0:hps_only_master_master_writedata
	wire  [31:0] hps_only_master_master_address;                                   // hps_only_master:master_address -> mm_interconnect_0:hps_only_master_master_address
	wire         hps_only_master_master_write;                                     // hps_only_master:master_write -> mm_interconnect_0:hps_only_master_master_write
	wire         hps_only_master_master_read;                                      // hps_only_master:master_read -> mm_interconnect_0:hps_only_master_master_read
	wire  [31:0] hps_only_master_master_readdata;                                  // mm_interconnect_0:hps_only_master_master_readdata -> hps_only_master:master_readdata
	wire   [3:0] hps_only_master_master_byteenable;                                // hps_only_master:master_byteenable -> mm_interconnect_0:hps_only_master_master_byteenable
	wire         hps_only_master_master_readdatavalid;                             // mm_interconnect_0:hps_only_master_master_readdatavalid -> hps_only_master:master_readdatavalid
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;                    // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;                     // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;                     // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;                    // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_arready;                    // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;                       // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rready;                     // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_bready;                     // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;                     // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;                     // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;                    // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire   [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;                     // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;                        // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;                      // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_awready;                    // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;                       // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;                     // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;                        // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;                     // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;                    // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;                      // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire   [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;                     // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire   [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;                     // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;                      // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;                     // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;                    // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire  [63:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;                      // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wready;                     // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire  [63:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;                      // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire  [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;                     // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;                    // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire   [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;                      // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire  [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;                     // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire   [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;                        // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;                     // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;                      // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_wlast;                      // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire         mm_interconnect_0_hps_0_f2h_axi_slave_rlast;                      // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire   [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;               // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;              // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_1_intr_capturer_0_avalon_slave_0_address;         // mm_interconnect_1:intr_capturer_0_avalon_slave_0_address -> intr_capturer_0:addr
	wire         mm_interconnect_1_intr_capturer_0_avalon_slave_0_read;            // mm_interconnect_1:intr_capturer_0_avalon_slave_0_read -> intr_capturer_0:read
	wire  [31:0] mm_interconnect_1_intr_capturer_0_avalon_slave_0_readdata;        // intr_capturer_0:rddata -> mm_interconnect_1:intr_capturer_0_avalon_slave_0_readdata
	wire         fpga_only_master_master_waitrequest;                              // mm_interconnect_1:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire  [31:0] fpga_only_master_master_writedata;                                // fpga_only_master:master_writedata -> mm_interconnect_1:fpga_only_master_master_writedata
	wire  [31:0] fpga_only_master_master_address;                                  // fpga_only_master:master_address -> mm_interconnect_1:fpga_only_master_master_address
	wire         fpga_only_master_master_write;                                    // fpga_only_master:master_write -> mm_interconnect_1:fpga_only_master_master_write
	wire         fpga_only_master_master_read;                                     // fpga_only_master:master_read -> mm_interconnect_1:fpga_only_master_master_read
	wire  [31:0] fpga_only_master_master_readdata;                                 // mm_interconnect_1:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire   [3:0] fpga_only_master_master_byteenable;                               // fpga_only_master:master_byteenable -> mm_interconnect_1:fpga_only_master_master_byteenable
	wire         fpga_only_master_master_readdatavalid;                            // mm_interconnect_1:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire  [31:0] mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_writedata;            // mm_interconnect_2:fifo_bridge_cpuM_cpus0_s0_writedata -> fifo_bridge_cpuM_cpus0:cpu1_writedata
	wire   [7:0] mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_address;              // mm_interconnect_2:fifo_bridge_cpuM_cpus0_s0_address -> fifo_bridge_cpuM_cpus0:cpu1_address
	wire         mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_write;                // mm_interconnect_2:fifo_bridge_cpuM_cpus0_s0_write -> fifo_bridge_cpuM_cpus0:cpu1_write
	wire         mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_read;                 // mm_interconnect_2:fifo_bridge_cpuM_cpus0_s0_read -> fifo_bridge_cpuM_cpus0:cpu1_read
	wire  [31:0] mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_readdata;             // fifo_bridge_cpuM_cpus0:cpu1_readdata -> mm_interconnect_2:fifo_bridge_cpuM_cpus0_s0_readdata
	wire         cpu_s0_data_master_waitrequest;                                   // mm_interconnect_2:cpu_s0_data_master_waitrequest -> cpu_s0:d_waitrequest
	wire  [31:0] cpu_s0_data_master_writedata;                                     // cpu_s0:d_writedata -> mm_interconnect_2:cpu_s0_data_master_writedata
	wire  [27:0] cpu_s0_data_master_address;                                       // cpu_s0:d_address -> mm_interconnect_2:cpu_s0_data_master_address
	wire         cpu_s0_data_master_write;                                         // cpu_s0:d_write -> mm_interconnect_2:cpu_s0_data_master_write
	wire         cpu_s0_data_master_read;                                          // cpu_s0:d_read -> mm_interconnect_2:cpu_s0_data_master_read
	wire  [31:0] cpu_s0_data_master_readdata;                                      // mm_interconnect_2:cpu_s0_data_master_readdata -> cpu_s0:d_readdata
	wire         cpu_s0_data_master_debugaccess;                                   // cpu_s0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_2:cpu_s0_data_master_debugaccess
	wire   [3:0] cpu_s0_data_master_byteenable;                                    // cpu_s0:d_byteenable -> mm_interconnect_2:cpu_s0_data_master_byteenable
	wire  [31:0] mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_writedata;           // mm_interconnect_2:fifo_bridge_cpus0_cpus1_s0_writedata -> fifo_bridge_cpus0_cpus1:cpu1_writedata
	wire   [7:0] mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_address;             // mm_interconnect_2:fifo_bridge_cpus0_cpus1_s0_address -> fifo_bridge_cpus0_cpus1:cpu1_address
	wire         mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_write;               // mm_interconnect_2:fifo_bridge_cpus0_cpus1_s0_write -> fifo_bridge_cpus0_cpus1:cpu1_write
	wire         mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_read;                // mm_interconnect_2:fifo_bridge_cpus0_cpus1_s0_read -> fifo_bridge_cpus0_cpus1:cpu1_read
	wire  [31:0] mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_readdata;            // fifo_bridge_cpus0_cpus1:cpu1_readdata -> mm_interconnect_2:fifo_bridge_cpus0_cpus1_s0_readdata
	wire         mm_interconnect_2_cpu_s0_jtag_debug_module_waitrequest;           // cpu_s0:jtag_debug_module_waitrequest -> mm_interconnect_2:cpu_s0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_2_cpu_s0_jtag_debug_module_writedata;             // mm_interconnect_2:cpu_s0_jtag_debug_module_writedata -> cpu_s0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_2_cpu_s0_jtag_debug_module_address;               // mm_interconnect_2:cpu_s0_jtag_debug_module_address -> cpu_s0:jtag_debug_module_address
	wire         mm_interconnect_2_cpu_s0_jtag_debug_module_write;                 // mm_interconnect_2:cpu_s0_jtag_debug_module_write -> cpu_s0:jtag_debug_module_write
	wire         mm_interconnect_2_cpu_s0_jtag_debug_module_read;                  // mm_interconnect_2:cpu_s0_jtag_debug_module_read -> cpu_s0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_2_cpu_s0_jtag_debug_module_readdata;              // cpu_s0:jtag_debug_module_readdata -> mm_interconnect_2:cpu_s0_jtag_debug_module_readdata
	wire         mm_interconnect_2_cpu_s0_jtag_debug_module_debugaccess;           // mm_interconnect_2:cpu_s0_jtag_debug_module_debugaccess -> cpu_s0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_2_cpu_s0_jtag_debug_module_byteenable;            // mm_interconnect_2:cpu_s0_jtag_debug_module_byteenable -> cpu_s0:jtag_debug_module_byteenable
	wire         mm_interconnect_2_s0_io_clockcrossing_bridge_s0_waitrequest;      // s0_io_clockCrossing_bridge:s0_waitrequest -> mm_interconnect_2:s0_io_clockCrossing_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_2_s0_io_clockcrossing_bridge_s0_burstcount;       // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_burstcount -> s0_io_clockCrossing_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_2_s0_io_clockcrossing_bridge_s0_writedata;        // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_writedata -> s0_io_clockCrossing_bridge:s0_writedata
	wire   [9:0] mm_interconnect_2_s0_io_clockcrossing_bridge_s0_address;          // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_address -> s0_io_clockCrossing_bridge:s0_address
	wire         mm_interconnect_2_s0_io_clockcrossing_bridge_s0_write;            // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_write -> s0_io_clockCrossing_bridge:s0_write
	wire         mm_interconnect_2_s0_io_clockcrossing_bridge_s0_read;             // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_read -> s0_io_clockCrossing_bridge:s0_read
	wire  [31:0] mm_interconnect_2_s0_io_clockcrossing_bridge_s0_readdata;         // s0_io_clockCrossing_bridge:s0_readdata -> mm_interconnect_2:s0_io_clockCrossing_bridge_s0_readdata
	wire         mm_interconnect_2_s0_io_clockcrossing_bridge_s0_debugaccess;      // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_debugaccess -> s0_io_clockCrossing_bridge:s0_debugaccess
	wire         mm_interconnect_2_s0_io_clockcrossing_bridge_s0_readdatavalid;    // s0_io_clockCrossing_bridge:s0_readdatavalid -> mm_interconnect_2:s0_io_clockCrossing_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_2_s0_io_clockcrossing_bridge_s0_byteenable;       // mm_interconnect_2:s0_io_clockCrossing_bridge_s0_byteenable -> s0_io_clockCrossing_bridge:s0_byteenable
	wire   [3:0] cpu_s0_instruction_master_burstcount;                             // cpu_s0:i_burstcount -> mm_interconnect_2:cpu_s0_instruction_master_burstcount
	wire         cpu_s0_instruction_master_waitrequest;                            // mm_interconnect_2:cpu_s0_instruction_master_waitrequest -> cpu_s0:i_waitrequest
	wire  [27:0] cpu_s0_instruction_master_address;                                // cpu_s0:i_address -> mm_interconnect_2:cpu_s0_instruction_master_address
	wire         cpu_s0_instruction_master_read;                                   // cpu_s0:i_read -> mm_interconnect_2:cpu_s0_instruction_master_read
	wire  [31:0] cpu_s0_instruction_master_readdata;                               // mm_interconnect_2:cpu_s0_instruction_master_readdata -> cpu_s0:i_readdata
	wire         cpu_s0_instruction_master_readdatavalid;                          // mm_interconnect_2:cpu_s0_instruction_master_readdatavalid -> cpu_s0:i_readdatavalid
	wire         mm_interconnect_2_sdram_clockcrossing_bridge_s0_waitrequest;      // sdram_clockCrossing_Bridge:s0_waitrequest -> mm_interconnect_2:sdram_clockCrossing_Bridge_s0_waitrequest
	wire   [3:0] mm_interconnect_2_sdram_clockcrossing_bridge_s0_burstcount;       // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_burstcount -> sdram_clockCrossing_Bridge:s0_burstcount
	wire  [31:0] mm_interconnect_2_sdram_clockcrossing_bridge_s0_writedata;        // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_writedata -> sdram_clockCrossing_Bridge:s0_writedata
	wire  [25:0] mm_interconnect_2_sdram_clockcrossing_bridge_s0_address;          // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_address -> sdram_clockCrossing_Bridge:s0_address
	wire         mm_interconnect_2_sdram_clockcrossing_bridge_s0_write;            // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_write -> sdram_clockCrossing_Bridge:s0_write
	wire         mm_interconnect_2_sdram_clockcrossing_bridge_s0_read;             // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_read -> sdram_clockCrossing_Bridge:s0_read
	wire  [31:0] mm_interconnect_2_sdram_clockcrossing_bridge_s0_readdata;         // sdram_clockCrossing_Bridge:s0_readdata -> mm_interconnect_2:sdram_clockCrossing_Bridge_s0_readdata
	wire         mm_interconnect_2_sdram_clockcrossing_bridge_s0_debugaccess;      // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_debugaccess -> sdram_clockCrossing_Bridge:s0_debugaccess
	wire         mm_interconnect_2_sdram_clockcrossing_bridge_s0_readdatavalid;    // sdram_clockCrossing_Bridge:s0_readdatavalid -> mm_interconnect_2:sdram_clockCrossing_Bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_2_sdram_clockcrossing_bridge_s0_byteenable;       // mm_interconnect_2:sdram_clockCrossing_Bridge_s0_byteenable -> sdram_clockCrossing_Bridge:s0_byteenable
	wire  [31:0] mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_writedata;            // mm_interconnect_3:fifo_bridge_cpuM_cpus0_s1_writedata -> fifo_bridge_cpuM_cpus0:cpu2_writedata
	wire   [7:0] mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_address;              // mm_interconnect_3:fifo_bridge_cpuM_cpus0_s1_address -> fifo_bridge_cpuM_cpus0:cpu2_address
	wire         mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_write;                // mm_interconnect_3:fifo_bridge_cpuM_cpus0_s1_write -> fifo_bridge_cpuM_cpus0:cpu2_write
	wire         mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_read;                 // mm_interconnect_3:fifo_bridge_cpuM_cpus0_s1_read -> fifo_bridge_cpuM_cpus0:cpu2_read
	wire  [31:0] mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_readdata;             // fifo_bridge_cpuM_cpus0:cpu2_readdata -> mm_interconnect_3:fifo_bridge_cpuM_cpus0_s1_readdata
	wire         hps_0_h2f_lw_axi_master_awvalid;                                  // hps_0:h2f_lw_AWVALID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awvalid
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                   // hps_0:h2f_lw_ARSIZE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arsize
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                   // hps_0:h2f_lw_ARLOCK -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arlock
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                  // hps_0:h2f_lw_AWCACHE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awcache
	wire         hps_0_h2f_lw_axi_master_arready;                                  // mm_interconnect_3:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                     // hps_0:h2f_lw_ARID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arid
	wire         hps_0_h2f_lw_axi_master_rready;                                   // hps_0:h2f_lw_RREADY -> mm_interconnect_3:hps_0_h2f_lw_axi_master_rready
	wire         hps_0_h2f_lw_axi_master_bready;                                   // hps_0:h2f_lw_BREADY -> mm_interconnect_3:hps_0_h2f_lw_axi_master_bready
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                   // hps_0:h2f_lw_AWSIZE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awsize
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                   // hps_0:h2f_lw_AWPROT -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awprot
	wire         hps_0_h2f_lw_axi_master_arvalid;                                  // hps_0:h2f_lw_ARVALID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arvalid
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                   // hps_0:h2f_lw_ARPROT -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arprot
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                      // mm_interconnect_3:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                    // hps_0:h2f_lw_ARLEN -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arlen
	wire         hps_0_h2f_lw_axi_master_awready;                                  // mm_interconnect_3:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                     // hps_0:h2f_lw_AWID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awid
	wire         hps_0_h2f_lw_axi_master_bvalid;                                   // mm_interconnect_3:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                      // hps_0:h2f_lw_WID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wid
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                   // hps_0:h2f_lw_AWLOCK -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                  // hps_0:h2f_lw_AWBURST -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awburst
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                    // mm_interconnect_3:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                    // hps_0:h2f_lw_WSTRB -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_rvalid;                                   // mm_interconnect_3:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                    // hps_0:h2f_lw_WDATA -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_wready;                                   // mm_interconnect_3:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                  // hps_0:h2f_lw_ARBURST -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arburst
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                    // mm_interconnect_3:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                   // hps_0:h2f_lw_ARADDR -> mm_interconnect_3:hps_0_h2f_lw_axi_master_araddr
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                  // hps_0:h2f_lw_ARCACHE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arcache
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                    // hps_0:h2f_lw_AWLEN -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awlen
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                   // hps_0:h2f_lw_AWADDR -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awaddr
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                      // mm_interconnect_3:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_wvalid;                                   // hps_0:h2f_lw_WVALID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wvalid
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                    // mm_interconnect_3:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire         hps_0_h2f_lw_axi_master_wlast;                                    // hps_0:h2f_lw_WLAST -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wlast
	wire         hps_0_h2f_lw_axi_master_rlast;                                    // mm_interconnect_3:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire  [31:0] mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_writedata;            // mm_interconnect_3:fifo_bridge_cpuM_cpus1_s1_writedata -> fifo_bridge_cpuM_cpus1:cpu2_writedata
	wire   [7:0] mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_address;              // mm_interconnect_3:fifo_bridge_cpuM_cpus1_s1_address -> fifo_bridge_cpuM_cpus1:cpu2_address
	wire         mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_write;                // mm_interconnect_3:fifo_bridge_cpuM_cpus1_s1_write -> fifo_bridge_cpuM_cpus1:cpu2_write
	wire         mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_read;                 // mm_interconnect_3:fifo_bridge_cpuM_cpus1_s1_read -> fifo_bridge_cpuM_cpus1:cpu2_read
	wire  [31:0] mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_readdata;             // fifo_bridge_cpuM_cpus1:cpu2_readdata -> mm_interconnect_3:fifo_bridge_cpuM_cpus1_s1_readdata
	wire  [31:0] mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_writedata;           // mm_interconnect_4:fifo_bridge_cpus0_cpus1_s1_writedata -> fifo_bridge_cpus0_cpus1:cpu2_writedata
	wire   [7:0] mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_address;             // mm_interconnect_4:fifo_bridge_cpus0_cpus1_s1_address -> fifo_bridge_cpus0_cpus1:cpu2_address
	wire         mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_write;               // mm_interconnect_4:fifo_bridge_cpus0_cpus1_s1_write -> fifo_bridge_cpus0_cpus1:cpu2_write
	wire         mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_read;                // mm_interconnect_4:fifo_bridge_cpus0_cpus1_s1_read -> fifo_bridge_cpus0_cpus1:cpu2_read
	wire  [31:0] mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_readdata;            // fifo_bridge_cpus0_cpus1:cpu2_readdata -> mm_interconnect_4:fifo_bridge_cpus0_cpus1_s1_readdata
	wire         cpu_s1_instruction_master_waitrequest;                            // mm_interconnect_4:cpu_s1_instruction_master_waitrequest -> cpu_s1:i_waitrequest
	wire  [27:0] cpu_s1_instruction_master_address;                                // cpu_s1:i_address -> mm_interconnect_4:cpu_s1_instruction_master_address
	wire         cpu_s1_instruction_master_read;                                   // cpu_s1:i_read -> mm_interconnect_4:cpu_s1_instruction_master_read
	wire  [31:0] cpu_s1_instruction_master_readdata;                               // mm_interconnect_4:cpu_s1_instruction_master_readdata -> cpu_s1:i_readdata
	wire         cpu_s1_instruction_master_readdatavalid;                          // mm_interconnect_4:cpu_s1_instruction_master_readdatavalid -> cpu_s1:i_readdatavalid
	wire  [31:0] mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_writedata;            // mm_interconnect_4:fifo_bridge_cpuM_cpus1_s0_writedata -> fifo_bridge_cpuM_cpus1:cpu1_writedata
	wire   [7:0] mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_address;              // mm_interconnect_4:fifo_bridge_cpuM_cpus1_s0_address -> fifo_bridge_cpuM_cpus1:cpu1_address
	wire         mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_write;                // mm_interconnect_4:fifo_bridge_cpuM_cpus1_s0_write -> fifo_bridge_cpuM_cpus1:cpu1_write
	wire         mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_read;                 // mm_interconnect_4:fifo_bridge_cpuM_cpus1_s0_read -> fifo_bridge_cpuM_cpus1:cpu1_read
	wire  [31:0] mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_readdata;             // fifo_bridge_cpuM_cpus1:cpu1_readdata -> mm_interconnect_4:fifo_bridge_cpuM_cpus1_s0_readdata
	wire         mm_interconnect_4_s1_io_clockcrossing_bridge_s0_waitrequest;      // s1_io_clockCrossing_bridge:s0_waitrequest -> mm_interconnect_4:s1_io_clockCrossing_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_4_s1_io_clockcrossing_bridge_s0_burstcount;       // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_burstcount -> s1_io_clockCrossing_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_4_s1_io_clockcrossing_bridge_s0_writedata;        // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_writedata -> s1_io_clockCrossing_bridge:s0_writedata
	wire   [9:0] mm_interconnect_4_s1_io_clockcrossing_bridge_s0_address;          // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_address -> s1_io_clockCrossing_bridge:s0_address
	wire         mm_interconnect_4_s1_io_clockcrossing_bridge_s0_write;            // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_write -> s1_io_clockCrossing_bridge:s0_write
	wire         mm_interconnect_4_s1_io_clockcrossing_bridge_s0_read;             // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_read -> s1_io_clockCrossing_bridge:s0_read
	wire  [31:0] mm_interconnect_4_s1_io_clockcrossing_bridge_s0_readdata;         // s1_io_clockCrossing_bridge:s0_readdata -> mm_interconnect_4:s1_io_clockCrossing_bridge_s0_readdata
	wire         mm_interconnect_4_s1_io_clockcrossing_bridge_s0_debugaccess;      // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_debugaccess -> s1_io_clockCrossing_bridge:s0_debugaccess
	wire         mm_interconnect_4_s1_io_clockcrossing_bridge_s0_readdatavalid;    // s1_io_clockCrossing_bridge:s0_readdatavalid -> mm_interconnect_4:s1_io_clockCrossing_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_4_s1_io_clockcrossing_bridge_s0_byteenable;       // mm_interconnect_4:s1_io_clockCrossing_bridge_s0_byteenable -> s1_io_clockCrossing_bridge:s0_byteenable
	wire  [31:0] mm_interconnect_4_onchip_sram_s1_writedata;                       // mm_interconnect_4:onchip_sram_s1_writedata -> onchip_sram:writedata
	wire  [16:0] mm_interconnect_4_onchip_sram_s1_address;                         // mm_interconnect_4:onchip_sram_s1_address -> onchip_sram:address
	wire         mm_interconnect_4_onchip_sram_s1_chipselect;                      // mm_interconnect_4:onchip_sram_s1_chipselect -> onchip_sram:chipselect
	wire         mm_interconnect_4_onchip_sram_s1_clken;                           // mm_interconnect_4:onchip_sram_s1_clken -> onchip_sram:clken
	wire         mm_interconnect_4_onchip_sram_s1_write;                           // mm_interconnect_4:onchip_sram_s1_write -> onchip_sram:write
	wire  [31:0] mm_interconnect_4_onchip_sram_s1_readdata;                        // onchip_sram:readdata -> mm_interconnect_4:onchip_sram_s1_readdata
	wire   [3:0] mm_interconnect_4_onchip_sram_s1_byteenable;                      // mm_interconnect_4:onchip_sram_s1_byteenable -> onchip_sram:byteenable
	wire         cpu_s1_data_master_waitrequest;                                   // mm_interconnect_4:cpu_s1_data_master_waitrequest -> cpu_s1:d_waitrequest
	wire  [31:0] cpu_s1_data_master_writedata;                                     // cpu_s1:d_writedata -> mm_interconnect_4:cpu_s1_data_master_writedata
	wire  [27:0] cpu_s1_data_master_address;                                       // cpu_s1:d_address -> mm_interconnect_4:cpu_s1_data_master_address
	wire         cpu_s1_data_master_write;                                         // cpu_s1:d_write -> mm_interconnect_4:cpu_s1_data_master_write
	wire         cpu_s1_data_master_read;                                          // cpu_s1:d_read -> mm_interconnect_4:cpu_s1_data_master_read
	wire  [31:0] cpu_s1_data_master_readdata;                                      // mm_interconnect_4:cpu_s1_data_master_readdata -> cpu_s1:d_readdata
	wire         cpu_s1_data_master_debugaccess;                                   // cpu_s1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_4:cpu_s1_data_master_debugaccess
	wire   [3:0] cpu_s1_data_master_byteenable;                                    // cpu_s1:d_byteenable -> mm_interconnect_4:cpu_s1_data_master_byteenable
	wire         mm_interconnect_4_cpu_s1_jtag_debug_module_waitrequest;           // cpu_s1:jtag_debug_module_waitrequest -> mm_interconnect_4:cpu_s1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_4_cpu_s1_jtag_debug_module_writedata;             // mm_interconnect_4:cpu_s1_jtag_debug_module_writedata -> cpu_s1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_4_cpu_s1_jtag_debug_module_address;               // mm_interconnect_4:cpu_s1_jtag_debug_module_address -> cpu_s1:jtag_debug_module_address
	wire         mm_interconnect_4_cpu_s1_jtag_debug_module_write;                 // mm_interconnect_4:cpu_s1_jtag_debug_module_write -> cpu_s1:jtag_debug_module_write
	wire         mm_interconnect_4_cpu_s1_jtag_debug_module_read;                  // mm_interconnect_4:cpu_s1_jtag_debug_module_read -> cpu_s1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_4_cpu_s1_jtag_debug_module_readdata;              // cpu_s1:jtag_debug_module_readdata -> mm_interconnect_4:cpu_s1_jtag_debug_module_readdata
	wire         mm_interconnect_4_cpu_s1_jtag_debug_module_debugaccess;           // mm_interconnect_4:cpu_s1_jtag_debug_module_debugaccess -> cpu_s1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_4_cpu_s1_jtag_debug_module_byteenable;            // mm_interconnect_4:cpu_s1_jtag_debug_module_byteenable -> cpu_s1:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_3_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_3_s0_writedata -> pwm_cpu_s0_3:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_3_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_3_s0_write -> pwm_cpu_s0_3:avs_s0_write
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_5_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_5_s0_writedata -> pwm_cpu_s0_5:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_5_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_5_s0_write -> pwm_cpu_s0_5:avs_s0_write
	wire   [0:0] s0_io_clockcrossing_bridge_m0_burstcount;                         // s0_io_clockCrossing_bridge:m0_burstcount -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_burstcount
	wire         s0_io_clockcrossing_bridge_m0_waitrequest;                        // mm_interconnect_5:s0_io_clockCrossing_bridge_m0_waitrequest -> s0_io_clockCrossing_bridge:m0_waitrequest
	wire   [9:0] s0_io_clockcrossing_bridge_m0_address;                            // s0_io_clockCrossing_bridge:m0_address -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_address
	wire  [31:0] s0_io_clockcrossing_bridge_m0_writedata;                          // s0_io_clockCrossing_bridge:m0_writedata -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_writedata
	wire         s0_io_clockcrossing_bridge_m0_write;                              // s0_io_clockCrossing_bridge:m0_write -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_write
	wire         s0_io_clockcrossing_bridge_m0_read;                               // s0_io_clockCrossing_bridge:m0_read -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_read
	wire  [31:0] s0_io_clockcrossing_bridge_m0_readdata;                           // mm_interconnect_5:s0_io_clockCrossing_bridge_m0_readdata -> s0_io_clockCrossing_bridge:m0_readdata
	wire         s0_io_clockcrossing_bridge_m0_debugaccess;                        // s0_io_clockCrossing_bridge:m0_debugaccess -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_debugaccess
	wire   [3:0] s0_io_clockcrossing_bridge_m0_byteenable;                         // s0_io_clockCrossing_bridge:m0_byteenable -> mm_interconnect_5:s0_io_clockCrossing_bridge_m0_byteenable
	wire         s0_io_clockcrossing_bridge_m0_readdatavalid;                      // mm_interconnect_5:s0_io_clockCrossing_bridge_m0_readdatavalid -> s0_io_clockCrossing_bridge:m0_readdatavalid
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_1_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_1_s0_writedata -> pwm_cpu_s0_1:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_1_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_1_s0_write -> pwm_cpu_s0_1:avs_s0_write
	wire  [31:0] mm_interconnect_5_pio_alivetest_cpu_s0_s1_writedata;              // mm_interconnect_5:pio_aliveTest_cpu_s0_s1_writedata -> pio_aliveTest_cpu_s0:writedata
	wire   [1:0] mm_interconnect_5_pio_alivetest_cpu_s0_s1_address;                // mm_interconnect_5:pio_aliveTest_cpu_s0_s1_address -> pio_aliveTest_cpu_s0:address
	wire         mm_interconnect_5_pio_alivetest_cpu_s0_s1_chipselect;             // mm_interconnect_5:pio_aliveTest_cpu_s0_s1_chipselect -> pio_aliveTest_cpu_s0:chipselect
	wire         mm_interconnect_5_pio_alivetest_cpu_s0_s1_write;                  // mm_interconnect_5:pio_aliveTest_cpu_s0_s1_write -> pio_aliveTest_cpu_s0:write_n
	wire  [31:0] mm_interconnect_5_pio_alivetest_cpu_s0_s1_readdata;               // pio_aliveTest_cpu_s0:readdata -> mm_interconnect_5:pio_aliveTest_cpu_s0_s1_readdata
	wire  [15:0] mm_interconnect_5_timer_cpu_s0_s1_writedata;                      // mm_interconnect_5:timer_cpu_s0_s1_writedata -> timer_cpu_s0:writedata
	wire   [2:0] mm_interconnect_5_timer_cpu_s0_s1_address;                        // mm_interconnect_5:timer_cpu_s0_s1_address -> timer_cpu_s0:address
	wire         mm_interconnect_5_timer_cpu_s0_s1_chipselect;                     // mm_interconnect_5:timer_cpu_s0_s1_chipselect -> timer_cpu_s0:chipselect
	wire         mm_interconnect_5_timer_cpu_s0_s1_write;                          // mm_interconnect_5:timer_cpu_s0_s1_write -> timer_cpu_s0:write_n
	wire  [15:0] mm_interconnect_5_timer_cpu_s0_s1_readdata;                       // timer_cpu_s0:readdata -> mm_interconnect_5:timer_cpu_s0_s1_readdata
	wire         mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_waitrequest; // jtag_uart_cpu_s0:av_waitrequest -> mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_writedata;   // mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_writedata -> jtag_uart_cpu_s0:av_writedata
	wire   [0:0] mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_address;     // mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_address -> jtag_uart_cpu_s0:av_address
	wire         mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_chipselect;  // mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_chipselect -> jtag_uart_cpu_s0:av_chipselect
	wire         mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_write;       // mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_write -> jtag_uart_cpu_s0:av_write_n
	wire         mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_read;        // mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_read -> jtag_uart_cpu_s0:av_read_n
	wire  [31:0] mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_readdata;    // jtag_uart_cpu_s0:av_readdata -> mm_interconnect_5:jtag_uart_cpu_s0_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_7_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_7_s0_writedata -> pwm_cpu_s0_7:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_7_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_7_s0_write -> pwm_cpu_s0_7:avs_s0_write
	wire         mm_interconnect_5_i2c_cpu_s0_mm_slave_waitrequest;                // i2c_cpu_s0:wb_ack_o -> mm_interconnect_5:i2c_cpu_s0_mm_slave_waitrequest
	wire   [7:0] mm_interconnect_5_i2c_cpu_s0_mm_slave_writedata;                  // mm_interconnect_5:i2c_cpu_s0_mm_slave_writedata -> i2c_cpu_s0:wb_dat_i
	wire   [2:0] mm_interconnect_5_i2c_cpu_s0_mm_slave_address;                    // mm_interconnect_5:i2c_cpu_s0_mm_slave_address -> i2c_cpu_s0:wb_adr_i
	wire         mm_interconnect_5_i2c_cpu_s0_mm_slave_chipselect;                 // mm_interconnect_5:i2c_cpu_s0_mm_slave_chipselect -> i2c_cpu_s0:wb_cyc_i
	wire         mm_interconnect_5_i2c_cpu_s0_mm_slave_write;                      // mm_interconnect_5:i2c_cpu_s0_mm_slave_write -> i2c_cpu_s0:wb_we_i
	wire   [7:0] mm_interconnect_5_i2c_cpu_s0_mm_slave_readdata;                   // i2c_cpu_s0:wb_dat_o -> mm_interconnect_5:i2c_cpu_s0_mm_slave_readdata
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_2_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_2_s0_writedata -> pwm_cpu_s0_2:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_2_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_2_s0_write -> pwm_cpu_s0_2:avs_s0_write
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_6_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_6_s0_writedata -> pwm_cpu_s0_6:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_6_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_6_s0_write -> pwm_cpu_s0_6:avs_s0_write
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_8_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_8_s0_writedata -> pwm_cpu_s0_8:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_8_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_8_s0_write -> pwm_cpu_s0_8:avs_s0_write
	wire  [31:0] mm_interconnect_5_pwm_cpu_s0_4_s0_writedata;                      // mm_interconnect_5:pwm_cpu_s0_4_s0_writedata -> pwm_cpu_s0_4:avs_s0_writedata
	wire         mm_interconnect_5_pwm_cpu_s0_4_s0_write;                          // mm_interconnect_5:pwm_cpu_s0_4_s0_write -> pwm_cpu_s0_4:avs_s0_write
	wire   [3:0] sdram_clockcrossing_bridge_m0_burstcount;                         // sdram_clockCrossing_Bridge:m0_burstcount -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_burstcount
	wire         sdram_clockcrossing_bridge_m0_waitrequest;                        // mm_interconnect_6:sdram_clockCrossing_Bridge_m0_waitrequest -> sdram_clockCrossing_Bridge:m0_waitrequest
	wire  [25:0] sdram_clockcrossing_bridge_m0_address;                            // sdram_clockCrossing_Bridge:m0_address -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_address
	wire  [31:0] sdram_clockcrossing_bridge_m0_writedata;                          // sdram_clockCrossing_Bridge:m0_writedata -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_writedata
	wire         sdram_clockcrossing_bridge_m0_write;                              // sdram_clockCrossing_Bridge:m0_write -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_write
	wire         sdram_clockcrossing_bridge_m0_read;                               // sdram_clockCrossing_Bridge:m0_read -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_read
	wire  [31:0] sdram_clockcrossing_bridge_m0_readdata;                           // mm_interconnect_6:sdram_clockCrossing_Bridge_m0_readdata -> sdram_clockCrossing_Bridge:m0_readdata
	wire         sdram_clockcrossing_bridge_m0_debugaccess;                        // sdram_clockCrossing_Bridge:m0_debugaccess -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_debugaccess
	wire   [3:0] sdram_clockcrossing_bridge_m0_byteenable;                         // sdram_clockCrossing_Bridge:m0_byteenable -> mm_interconnect_6:sdram_clockCrossing_Bridge_m0_byteenable
	wire         sdram_clockcrossing_bridge_m0_readdatavalid;                      // mm_interconnect_6:sdram_clockCrossing_Bridge_m0_readdatavalid -> sdram_clockCrossing_Bridge:m0_readdatavalid
	wire         mm_interconnect_6_sdram_s1_waitrequest;                           // sdram:za_waitrequest -> mm_interconnect_6:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_6_sdram_s1_writedata;                             // mm_interconnect_6:sdram_s1_writedata -> sdram:az_data
	wire  [24:0] mm_interconnect_6_sdram_s1_address;                               // mm_interconnect_6:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_6_sdram_s1_chipselect;                            // mm_interconnect_6:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_6_sdram_s1_write;                                 // mm_interconnect_6:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_6_sdram_s1_read;                                  // mm_interconnect_6:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_6_sdram_s1_readdata;                              // sdram:za_data -> mm_interconnect_6:sdram_s1_readdata
	wire         mm_interconnect_6_sdram_s1_readdatavalid;                         // sdram:za_valid -> mm_interconnect_6:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_6_sdram_s1_byteenable;                            // mm_interconnect_6:sdram_s1_byteenable -> sdram:az_be_n
	wire   [0:0] s1_io_clockcrossing_bridge_m0_burstcount;                         // s1_io_clockCrossing_bridge:m0_burstcount -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_burstcount
	wire         s1_io_clockcrossing_bridge_m0_waitrequest;                        // mm_interconnect_7:s1_io_clockCrossing_bridge_m0_waitrequest -> s1_io_clockCrossing_bridge:m0_waitrequest
	wire   [9:0] s1_io_clockcrossing_bridge_m0_address;                            // s1_io_clockCrossing_bridge:m0_address -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_address
	wire  [31:0] s1_io_clockcrossing_bridge_m0_writedata;                          // s1_io_clockCrossing_bridge:m0_writedata -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_writedata
	wire         s1_io_clockcrossing_bridge_m0_write;                              // s1_io_clockCrossing_bridge:m0_write -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_write
	wire         s1_io_clockcrossing_bridge_m0_read;                               // s1_io_clockCrossing_bridge:m0_read -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_read
	wire  [31:0] s1_io_clockcrossing_bridge_m0_readdata;                           // mm_interconnect_7:s1_io_clockCrossing_bridge_m0_readdata -> s1_io_clockCrossing_bridge:m0_readdata
	wire         s1_io_clockcrossing_bridge_m0_debugaccess;                        // s1_io_clockCrossing_bridge:m0_debugaccess -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_debugaccess
	wire   [3:0] s1_io_clockcrossing_bridge_m0_byteenable;                         // s1_io_clockCrossing_bridge:m0_byteenable -> mm_interconnect_7:s1_io_clockCrossing_bridge_m0_byteenable
	wire         s1_io_clockcrossing_bridge_m0_readdatavalid;                      // mm_interconnect_7:s1_io_clockCrossing_bridge_m0_readdatavalid -> s1_io_clockCrossing_bridge:m0_readdatavalid
	wire         mm_interconnect_7_i2c_cpu_s1_mm_slave_waitrequest;                // i2c_cpu_s1:wb_ack_o -> mm_interconnect_7:i2c_cpu_s1_mm_slave_waitrequest
	wire   [7:0] mm_interconnect_7_i2c_cpu_s1_mm_slave_writedata;                  // mm_interconnect_7:i2c_cpu_s1_mm_slave_writedata -> i2c_cpu_s1:wb_dat_i
	wire   [2:0] mm_interconnect_7_i2c_cpu_s1_mm_slave_address;                    // mm_interconnect_7:i2c_cpu_s1_mm_slave_address -> i2c_cpu_s1:wb_adr_i
	wire         mm_interconnect_7_i2c_cpu_s1_mm_slave_chipselect;                 // mm_interconnect_7:i2c_cpu_s1_mm_slave_chipselect -> i2c_cpu_s1:wb_cyc_i
	wire         mm_interconnect_7_i2c_cpu_s1_mm_slave_write;                      // mm_interconnect_7:i2c_cpu_s1_mm_slave_write -> i2c_cpu_s1:wb_we_i
	wire   [7:0] mm_interconnect_7_i2c_cpu_s1_mm_slave_readdata;                   // i2c_cpu_s1:wb_dat_o -> mm_interconnect_7:i2c_cpu_s1_mm_slave_readdata
	wire  [15:0] mm_interconnect_7_timer_cpu_s1_s1_writedata;                      // mm_interconnect_7:timer_cpu_s1_s1_writedata -> timer_cpu_s1:writedata
	wire   [2:0] mm_interconnect_7_timer_cpu_s1_s1_address;                        // mm_interconnect_7:timer_cpu_s1_s1_address -> timer_cpu_s1:address
	wire         mm_interconnect_7_timer_cpu_s1_s1_chipselect;                     // mm_interconnect_7:timer_cpu_s1_s1_chipselect -> timer_cpu_s1:chipselect
	wire         mm_interconnect_7_timer_cpu_s1_s1_write;                          // mm_interconnect_7:timer_cpu_s1_s1_write -> timer_cpu_s1:write_n
	wire  [15:0] mm_interconnect_7_timer_cpu_s1_s1_readdata;                       // timer_cpu_s1:readdata -> mm_interconnect_7:timer_cpu_s1_s1_readdata
	wire         mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_waitrequest; // jtag_uart_cpu_s1:av_waitrequest -> mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_writedata;   // mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_writedata -> jtag_uart_cpu_s1:av_writedata
	wire   [0:0] mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_address;     // mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_address -> jtag_uart_cpu_s1:av_address
	wire         mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_chipselect;  // mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_chipselect -> jtag_uart_cpu_s1:av_chipselect
	wire         mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_write;       // mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_write -> jtag_uart_cpu_s1:av_write_n
	wire         mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_read;        // mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_read -> jtag_uart_cpu_s1:av_read_n
	wire  [31:0] mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_readdata;    // jtag_uart_cpu_s1:av_readdata -> mm_interconnect_7:jtag_uart_cpu_s1_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_7_pio_alivetest_cpu_s1_s1_writedata;              // mm_interconnect_7:pio_aliveTest_cpu_s1_s1_writedata -> pio_aliveTest_cpu_s1:writedata
	wire   [1:0] mm_interconnect_7_pio_alivetest_cpu_s1_s1_address;                // mm_interconnect_7:pio_aliveTest_cpu_s1_s1_address -> pio_aliveTest_cpu_s1:address
	wire         mm_interconnect_7_pio_alivetest_cpu_s1_s1_chipselect;             // mm_interconnect_7:pio_aliveTest_cpu_s1_s1_chipselect -> pio_aliveTest_cpu_s1:chipselect
	wire         mm_interconnect_7_pio_alivetest_cpu_s1_s1_write;                  // mm_interconnect_7:pio_aliveTest_cpu_s1_s1_write -> pio_aliveTest_cpu_s1:write_n
	wire  [31:0] mm_interconnect_7_pio_alivetest_cpu_s1_s1_readdata;               // pio_aliveTest_cpu_s1:readdata -> mm_interconnect_7:pio_aliveTest_cpu_s1_s1_readdata
	wire  [31:0] hps_0_f2h_irq0_irq;                                               // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                               // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire  [31:0] intr_capturer_0_interrupt_receiver_irq;                           // irq_mapper_002:sender_irq -> intr_capturer_0:interrupt_in
	wire         irq_mapper_003_receiver2_irq;                                     // fifo_bridge_cpuM_cpus0:cpu1_irq -> irq_mapper_003:receiver2_irq
	wire         irq_mapper_003_receiver3_irq;                                     // fifo_bridge_cpus0_cpus1:cpu1_irq -> irq_mapper_003:receiver3_irq
	wire  [31:0] cpu_s0_d_irq_irq;                                                 // irq_mapper_003:sender_irq -> cpu_s0:d_irq
	wire         irq_mapper_004_receiver2_irq;                                     // fifo_bridge_cpuM_cpus1:cpu1_irq -> irq_mapper_004:receiver2_irq
	wire         irq_mapper_004_receiver3_irq;                                     // fifo_bridge_cpus0_cpus1:cpu2_irq -> irq_mapper_004:receiver3_irq
	wire  [31:0] cpu_s1_d_irq_irq;                                                 // irq_mapper_004:sender_irq -> cpu_s1:d_irq
	wire         irq_mapper_003_receiver0_irq;                                     // irq_synchronizer:sender_irq -> irq_mapper_003:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                    // timer_cpu_s0:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_003_receiver1_irq;                                     // irq_synchronizer_001:sender_irq -> irq_mapper_003:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                // jtag_uart_cpu_s0:av_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_003_receiver4_irq;                                     // irq_synchronizer_002:sender_irq -> irq_mapper_003:receiver4_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                // i2c_cpu_s0:wb_inta_o -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_004_receiver0_irq;                                     // irq_synchronizer_003:sender_irq -> irq_mapper_004:receiver0_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                // timer_cpu_s1:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_004_receiver1_irq;                                     // irq_synchronizer_004:sender_irq -> irq_mapper_004:receiver1_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                // jtag_uart_cpu_s1:av_irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_004_receiver4_irq;                                     // irq_synchronizer_005:sender_irq -> irq_mapper_004:receiver4_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                                // i2c_cpu_s1:wb_inta_o -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver0_irq;                                         // fifo_bridge_cpuM_cpus0:cpu2_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver1_irq]
	wire         irq_mapper_receiver1_irq;                                         // fifo_bridge_cpuM_cpus1:cpu2_irq -> [irq_mapper:receiver1_irq, irq_mapper_002:receiver0_irq]
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [cpu_s0:reset_n, cpu_s1:reset_n, fifo_bridge_cpuM_cpus0:reset, fifo_bridge_cpuM_cpus1:reset, fifo_bridge_cpus0_cpus1:reset, intr_capturer_0:rst_n, irq_mapper_002:reset, irq_mapper_003:reset, irq_mapper_004:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, mm_interconnect_0:hps_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:hps_only_master_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:intr_capturer_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:cpu_s0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_3:fifo_bridge_cpuM_cpus0_clock_reset_reset_bridge_in_reset_reset, mm_interconnect_4:cpu_s1_reset_n_reset_bridge_in_reset_reset, onchip_sram:reset, rst_translator:in_reset, s0_io_clockCrossing_bridge:s0_reset, s1_io_clockCrossing_bridge:s0_reset, sdram_clockCrossing_Bridge:s0_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [cpu_s0:reset_req, cpu_s1:reset_req, onchip_sram:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [i2c_cpu_s0:wb_rst_i, i2c_cpu_s1:wb_rst_i, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, jtag_uart_cpu_s0:rst_n, jtag_uart_cpu_s1:rst_n, mm_interconnect_5:s0_io_clockCrossing_bridge_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_7:s1_io_clockCrossing_bridge_m0_reset_reset_bridge_in_reset_reset, pio_aliveTest_cpu_s0:reset_n, pio_aliveTest_cpu_s1:reset_n, s0_io_clockCrossing_bridge:m0_reset, s1_io_clockCrossing_bridge:m0_reset, timer_cpu_s0:reset_n, timer_cpu_s1:reset_n]
	wire         rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> [mm_interconnect_6:sdram_clockCrossing_Bridge_m0_reset_reset_bridge_in_reset_reset, sdram:reset_n, sdram_clockCrossing_Bridge:m0_reset]
	wire         rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> [pwm_pll:rst, sdram_pll:rst, system_pll:rst]
	wire         rst_controller_004_reset_out_reset;                               // rst_controller_004:reset_out -> [mm_interconnect_5:pwm_cpu_s0_1_clock_reset_reset_bridge_in_reset_reset, pwm_cpu_s0_1:reset, pwm_cpu_s0_2:reset, pwm_cpu_s0_3:reset, pwm_cpu_s0_4:reset, pwm_cpu_s0_5:reset, pwm_cpu_s0_6:reset, pwm_cpu_s0_7:reset, pwm_cpu_s0_8:reset]
	wire         rst_controller_005_reset_out_reset;                               // rst_controller_005:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_3:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),              //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),             // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),              //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),          //   f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                                  //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),         //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),           //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),           //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),           //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),           //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),           //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),           //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),            //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),         //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),         //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),         //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),           //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),           //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),           //                    .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),             //                    .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),             //                    .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),             //                    .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),             //                    .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),             //                    .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),             //                    .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),             //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),              //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),              //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),             //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),              //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),              //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),              //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),              //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),              //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),              //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),              //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),              //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),              //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),              //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),             //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),             //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),             //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),             //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),            //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),           //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),           //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),            //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),             //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),             //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),             //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),             //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),             //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),             //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),          //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),          //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),          //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),          //                    .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),          //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),          //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),          //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //           h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                                       //       h2f_axi_clock.clk
		.h2f_AWID                 (),                                              //      h2f_axi_master.awid
		.h2f_AWADDR               (),                                              //                    .awaddr
		.h2f_AWLEN                (),                                              //                    .awlen
		.h2f_AWSIZE               (),                                              //                    .awsize
		.h2f_AWBURST              (),                                              //                    .awburst
		.h2f_AWLOCK               (),                                              //                    .awlock
		.h2f_AWCACHE              (),                                              //                    .awcache
		.h2f_AWPROT               (),                                              //                    .awprot
		.h2f_AWVALID              (),                                              //                    .awvalid
		.h2f_AWREADY              (),                                              //                    .awready
		.h2f_WID                  (),                                              //                    .wid
		.h2f_WDATA                (),                                              //                    .wdata
		.h2f_WSTRB                (),                                              //                    .wstrb
		.h2f_WLAST                (),                                              //                    .wlast
		.h2f_WVALID               (),                                              //                    .wvalid
		.h2f_WREADY               (),                                              //                    .wready
		.h2f_BID                  (),                                              //                    .bid
		.h2f_BRESP                (),                                              //                    .bresp
		.h2f_BVALID               (),                                              //                    .bvalid
		.h2f_BREADY               (),                                              //                    .bready
		.h2f_ARID                 (),                                              //                    .arid
		.h2f_ARADDR               (),                                              //                    .araddr
		.h2f_ARLEN                (),                                              //                    .arlen
		.h2f_ARSIZE               (),                                              //                    .arsize
		.h2f_ARBURST              (),                                              //                    .arburst
		.h2f_ARLOCK               (),                                              //                    .arlock
		.h2f_ARCACHE              (),                                              //                    .arcache
		.h2f_ARPROT               (),                                              //                    .arprot
		.h2f_ARVALID              (),                                              //                    .arvalid
		.h2f_ARREADY              (),                                              //                    .arready
		.h2f_RID                  (),                                              //                    .rid
		.h2f_RDATA                (),                                              //                    .rdata
		.h2f_RRESP                (),                                              //                    .rresp
		.h2f_RLAST                (),                                              //                    .rlast
		.h2f_RVALID               (),                                              //                    .rvalid
		.h2f_RREADY               (),                                              //                    .rready
		.f2h_axi_clk              (clk_clk),                                       //       f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //       f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                    .awaddr
		.f2h_AWLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                    .awlen
		.f2h_AWSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                    .awsize
		.f2h_AWBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                    .awburst
		.f2h_AWLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                    .awlock
		.f2h_AWCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                    .awcache
		.f2h_AWPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                    .awprot
		.f2h_AWVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                    .awvalid
		.f2h_AWREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                    .awready
		.f2h_AWUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                    .awuser
		.f2h_WID                  (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                    .wid
		.f2h_WDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                    .wdata
		.f2h_WSTRB                (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                    .wstrb
		.f2h_WLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                    .wlast
		.f2h_WVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                    .wvalid
		.f2h_WREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                    .wready
		.f2h_BID                  (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                    .bid
		.f2h_BRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                    .bresp
		.f2h_BVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                    .bvalid
		.f2h_BREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                    .bready
		.f2h_ARID                 (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                    .arid
		.f2h_ARADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                    .araddr
		.f2h_ARLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                    .arlen
		.f2h_ARSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                    .arsize
		.f2h_ARBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                    .arburst
		.f2h_ARLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                    .arlock
		.f2h_ARCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                    .arcache
		.f2h_ARPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                    .arprot
		.f2h_ARVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                    .arvalid
		.f2h_ARREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                    .arready
		.f2h_ARUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                    .aruser
		.f2h_RID                  (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                    .rid
		.f2h_RDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                    .rdata
		.f2h_RRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                    .rresp
		.f2h_RLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                    .rlast
		.f2h_RVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                    .rvalid
		.f2h_RREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                                       //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                            //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                             //            f2h_irq1.irq
	);

	soc_system_onchip_sram onchip_sram (
		.clk        (system_pll_outclk0_clk),                      //   clk1.clk
		.address    (mm_interconnect_4_onchip_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_4_onchip_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_4_onchip_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_4_onchip_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_4_onchip_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_4_onchip_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_4_onchip_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)           //       .reset_req
	);

	soc_system_hps_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) hps_only_master (
		.clk_clk              (system_pll_outclk0_clk),               //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                       //    clk_reset.reset
		.master_address       (hps_only_master_master_address),       //       master.address
		.master_readdata      (hps_only_master_master_readdata),      //             .readdata
		.master_read          (hps_only_master_master_read),          //             .read
		.master_write         (hps_only_master_master_write),         //             .write
		.master_writedata     (hps_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (hps_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (hps_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (hps_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                      // master_reset.reset
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (system_pll_outclk0_clk),                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_hps_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (system_pll_outclk0_clk),                //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                        //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	intr_capturer #(
		.NUM_INTR (32)
	) intr_capturer_0 (
		.clk          (system_pll_outclk0_clk),                                    //              clock.clk
		.rst_n        (~rst_controller_reset_out_reset),                           //         reset_sink.reset_n
		.addr         (mm_interconnect_1_intr_capturer_0_avalon_slave_0_address),  //     avalon_slave_0.address
		.read         (mm_interconnect_1_intr_capturer_0_avalon_slave_0_read),     //                   .read
		.rddata       (mm_interconnect_1_intr_capturer_0_avalon_slave_0_readdata), //                   .readdata
		.interrupt_in (intr_capturer_0_interrupt_receiver_irq)                     // interrupt_receiver.irq
	);

	soc_system_pio_aliveTest_cpu_s0 pio_alivetest_cpu_s0 (
		.clk        (system_pll_outclk1_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_5_pio_alivetest_cpu_s0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_5_pio_alivetest_cpu_s0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_5_pio_alivetest_cpu_s0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_5_pio_alivetest_cpu_s0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_5_pio_alivetest_cpu_s0_s1_readdata),   //                    .readdata
		.out_port   (pio_alivetest_cpu_s0_extcon_export)                    // external_connection.export
	);

	soc_system_cpu_s0 cpu_s0 (
		.clk                                   (system_pll_outclk0_clk),                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_s0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_s0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_s0_data_master_read),                                //                          .read
		.d_readdata                            (cpu_s0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_s0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_s0_data_master_write),                               //                          .write
		.d_writedata                           (cpu_s0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_s0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_s0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_s0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_s0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_s0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_burstcount                          (cpu_s0_instruction_master_burstcount),                   //                          .burstcount
		.i_readdatavalid                       (cpu_s0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_s0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                       //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_2_cpu_s0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_2_cpu_s0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_2_cpu_s0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_2_cpu_s0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_2_cpu_s0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_2_cpu_s0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_2_cpu_s0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_2_cpu_s0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	soc_system_timer_cpu_s0 timer_cpu_s0 (
		.clk        (system_pll_outclk1_clk),                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_5_timer_cpu_s0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_5_timer_cpu_s0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_5_timer_cpu_s0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_5_timer_cpu_s0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_5_timer_cpu_s0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                 //   irq.irq
	);

	soc_system_jtag_uart_cpu_s0 jtag_uart_cpu_s0 (
		.clk            (system_pll_outclk1_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                                 //               irq.irq
	);

	soc_system_sdram sdram (
		.clk            (sdram_pll_outclk0_clk),                    //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_6_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_6_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_6_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_6_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_6_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_6_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_6_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_6_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_6_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	CPU_FiFo_Bridge fifo_bridge_cpum_cpus0 (
		.clk            (system_pll_outclk0_clk),                                //       clock.clk
		.reset          (rst_controller_reset_out_reset),                        // clock_reset.reset
		.cpu1_address   (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_address),   //          s0.address
		.cpu1_read      (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_read),      //            .read
		.cpu1_readdata  (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_readdata),  //            .readdata
		.cpu1_write     (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_write),     //            .write
		.cpu1_writedata (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_writedata), //            .writedata
		.cpu1_irq       (irq_mapper_003_receiver2_irq),                          //        irq0.irq
		.cpu2_address   (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_address),   //          s1.address
		.cpu2_read      (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_read),      //            .read
		.cpu2_readdata  (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_readdata),  //            .readdata
		.cpu2_writedata (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_writedata), //            .writedata
		.cpu2_write     (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_write),     //            .write
		.cpu2_irq       (irq_mapper_receiver0_irq)                               //        irq1.irq
	);

	soc_system_cpu_s1 cpu_s1 (
		.clk                                   (system_pll_outclk0_clk),                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_s1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_s1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_s1_data_master_read),                                //                          .read
		.d_readdata                            (cpu_s1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_s1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_s1_data_master_write),                               //                          .write
		.d_writedata                           (cpu_s1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_s1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_s1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_s1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_s1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_s1_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_s1_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_s1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                       //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_4_cpu_s1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_4_cpu_s1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_4_cpu_s1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_4_cpu_s1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_4_cpu_s1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_4_cpu_s1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_4_cpu_s1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_4_cpu_s1_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	soc_system_timer_cpu_s0 timer_cpu_s1 (
		.clk        (system_pll_outclk1_clk),                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_7_timer_cpu_s1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_7_timer_cpu_s1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_7_timer_cpu_s1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_7_timer_cpu_s1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_7_timer_cpu_s1_s1_write),     //      .write_n
		.irq        (irq_synchronizer_003_receiver_irq)             //   irq.irq
	);

	soc_system_jtag_uart_cpu_s0 jtag_uart_cpu_s1 (
		.clk            (system_pll_outclk1_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_004_receiver_irq)                                 //               irq.irq
	);

	soc_system_pio_aliveTest_cpu_s0 pio_alivetest_cpu_s1 (
		.clk        (system_pll_outclk1_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_7_pio_alivetest_cpu_s1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_7_pio_alivetest_cpu_s1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_7_pio_alivetest_cpu_s1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_7_pio_alivetest_cpu_s1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_7_pio_alivetest_cpu_s1_s1_readdata),   //                    .readdata
		.out_port   (pio_alivetest_cpu_s1_extcon_export)                    // external_connection.export
	);

	CPU_FiFo_Bridge fifo_bridge_cpus0_cpus1 (
		.clk            (system_pll_outclk0_clk),                                 //       clock.clk
		.reset          (rst_controller_reset_out_reset),                         // clock_reset.reset
		.cpu1_address   (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_address),   //          s0.address
		.cpu1_read      (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_read),      //            .read
		.cpu1_readdata  (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_readdata),  //            .readdata
		.cpu1_write     (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_write),     //            .write
		.cpu1_writedata (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_writedata), //            .writedata
		.cpu1_irq       (irq_mapper_003_receiver3_irq),                           //        irq0.irq
		.cpu2_address   (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_address),   //          s1.address
		.cpu2_read      (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_read),      //            .read
		.cpu2_readdata  (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_readdata),  //            .readdata
		.cpu2_writedata (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_writedata), //            .writedata
		.cpu2_write     (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_write),     //            .write
		.cpu2_irq       (irq_mapper_004_receiver3_irq)                            //        irq1.irq
	);

	CPU_FiFo_Bridge fifo_bridge_cpum_cpus1 (
		.clk            (system_pll_outclk0_clk),                                //       clock.clk
		.reset          (rst_controller_reset_out_reset),                        // clock_reset.reset
		.cpu1_address   (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_address),   //          s0.address
		.cpu1_read      (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_read),      //            .read
		.cpu1_readdata  (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_readdata),  //            .readdata
		.cpu1_write     (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_write),     //            .write
		.cpu1_writedata (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_writedata), //            .writedata
		.cpu1_irq       (irq_mapper_004_receiver2_irq),                          //        irq0.irq
		.cpu2_address   (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_address),   //          s1.address
		.cpu2_read      (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_read),      //            .read
		.cpu2_readdata  (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_readdata),  //            .readdata
		.cpu2_writedata (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_writedata), //            .writedata
		.cpu2_write     (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_write),     //            .write
		.cpu2_irq       (irq_mapper_receiver1_irq)                               //        irq1.irq
	);

	soc_system_system_pll system_pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (system_pll_outclk0_clk),             // outclk0.clk
		.outclk_1 (system_pll_outclk1_clk),             // outclk1.clk
		.locked   (system_pll_locked_export)            //  locked.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) s0_io_clockcrossing_bridge (
		.m0_clk           (system_pll_outclk1_clk),                                        //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (system_pll_outclk0_clk),                                        //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (s0_io_clockcrossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (s0_io_clockcrossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (s0_io_clockcrossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (s0_io_clockcrossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (s0_io_clockcrossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (s0_io_clockcrossing_bridge_m0_address),                         //         .address
		.m0_write         (s0_io_clockcrossing_bridge_m0_write),                           //         .write
		.m0_read          (s0_io_clockcrossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (s0_io_clockcrossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (s0_io_clockcrossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (26),
		.BURSTCOUNT_WIDTH    (4),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (16),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) sdram_clockcrossing_bridge (
		.m0_clk           (sdram_pll_outclk0_clk),                                         //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (system_pll_outclk0_clk),                                        //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_2_sdram_clockcrossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_2_sdram_clockcrossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_2_sdram_clockcrossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_2_sdram_clockcrossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_2_sdram_clockcrossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_2_sdram_clockcrossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_2_sdram_clockcrossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_2_sdram_clockcrossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_2_sdram_clockcrossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_2_sdram_clockcrossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (sdram_clockcrossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (sdram_clockcrossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (sdram_clockcrossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (sdram_clockcrossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (sdram_clockcrossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (sdram_clockcrossing_bridge_m0_address),                         //         .address
		.m0_write         (sdram_clockcrossing_bridge_m0_write),                           //         .write
		.m0_read          (sdram_clockcrossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (sdram_clockcrossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (sdram_clockcrossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	soc_system_sdram_pll sdram_pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (sdram_pll_outclk0_clk),              // outclk0.clk
		.outclk_1 (clk_sdram_clk),                      // outclk1.clk
		.locked   (sdram_pll_locked_export)             //  locked.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) s1_io_clockcrossing_bridge (
		.m0_clk           (system_pll_outclk1_clk),                                        //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (system_pll_outclk0_clk),                                        //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (s1_io_clockcrossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (s1_io_clockcrossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (s1_io_clockcrossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (s1_io_clockcrossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (s1_io_clockcrossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (s1_io_clockcrossing_bridge_m0_address),                         //         .address
		.m0_write         (s1_io_clockcrossing_bridge_m0_write),                           //         .write
		.m0_read          (s1_io_clockcrossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (s1_io_clockcrossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (s1_io_clockcrossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	oc_i2c_master i2c_cpu_s0 (
		.wb_clk_i  (system_pll_outclk1_clk),                            //           mm_clk.clk
		.wb_rst_i  (rst_controller_001_reset_out_reset),                //     mm_clk_reset.reset
		.wb_dat_i  (mm_interconnect_5_i2c_cpu_s0_mm_slave_writedata),   //         mm_slave.writedata
		.wb_dat_o  (mm_interconnect_5_i2c_cpu_s0_mm_slave_readdata),    //                 .readdata
		.wb_we_i   (mm_interconnect_5_i2c_cpu_s0_mm_slave_write),       //                 .write
		.wb_cyc_i  (mm_interconnect_5_i2c_cpu_s0_mm_slave_chipselect),  //                 .chipselect
		.wb_ack_o  (mm_interconnect_5_i2c_cpu_s0_mm_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i  (mm_interconnect_5_i2c_cpu_s0_mm_slave_address),     //                 .address
		.scl       (i2c_cpu_s0_i2c_exports_scl),                        //      i2c_exports.export
		.sda       (i2c_cpu_s0_i2c_exports_sda),                        //                 .export
		.wb_inta_o (irq_synchronizer_002_receiver_irq)                  // interrupt_sender.irq
	);

	oc_i2c_master i2c_cpu_s1 (
		.wb_clk_i  (system_pll_outclk1_clk),                            //           mm_clk.clk
		.wb_rst_i  (rst_controller_001_reset_out_reset),                //     mm_clk_reset.reset
		.wb_dat_i  (mm_interconnect_7_i2c_cpu_s1_mm_slave_writedata),   //         mm_slave.writedata
		.wb_dat_o  (mm_interconnect_7_i2c_cpu_s1_mm_slave_readdata),    //                 .readdata
		.wb_we_i   (mm_interconnect_7_i2c_cpu_s1_mm_slave_write),       //                 .write
		.wb_cyc_i  (mm_interconnect_7_i2c_cpu_s1_mm_slave_chipselect),  //                 .chipselect
		.wb_ack_o  (mm_interconnect_7_i2c_cpu_s1_mm_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i  (mm_interconnect_7_i2c_cpu_s1_mm_slave_address),     //                 .address
		.scl       (i2c_cpu_s1_i2c_exports_scl),                        //      i2c_exports.export
		.sda       (i2c_cpu_s1_i2c_exports_sda),                        //                 .export
		.wb_inta_o (irq_synchronizer_005_receiver_irq)                  // interrupt_sender.irq
	);

	pwm pwm_cpu_s0_1 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_1_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_1_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_1_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	soc_system_pwm_pll pwm_pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (pwm_pll_outclk0_clk),                // outclk0.clk
		.locked   ()                                    //  locked.export
	);

	pwm pwm_cpu_s0_2 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_2_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_2_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_2_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	pwm pwm_cpu_s0_3 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_3_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_3_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_3_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	pwm pwm_cpu_s0_4 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_4_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_4_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_4_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	pwm pwm_cpu_s0_5 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_5_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_5_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_5_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	pwm pwm_cpu_s0_6 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_6_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_6_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_6_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	pwm pwm_cpu_s0_7 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_7_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_7_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_7_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	pwm pwm_cpu_s0_8 (
		.clk              (pwm_pll_outclk0_clk),                         //       clock.clk
		.reset            (rst_controller_004_reset_out_reset),          // clock_reset.reset
		.avs_s0_write     (mm_interconnect_5_pwm_cpu_s0_8_s0_write),     //          s0.write
		.avs_s0_writedata (mm_interconnect_5_pwm_cpu_s0_8_s0_writedata), //            .writedata
		.out_signal       (pwm_cpu_s0_8_conduit_end_readdatavalid_n)     // conduit_end.readdatavalid_n
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                                            (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                                           hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                          (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                                              .awaddr
		.hps_0_f2h_axi_slave_awlen                                           (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                                              .awlen
		.hps_0_f2h_axi_slave_awsize                                          (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                                              .awsize
		.hps_0_f2h_axi_slave_awburst                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                                              .awburst
		.hps_0_f2h_axi_slave_awlock                                          (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                                              .awlock
		.hps_0_f2h_axi_slave_awcache                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                                              .awcache
		.hps_0_f2h_axi_slave_awprot                                          (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                                              .awprot
		.hps_0_f2h_axi_slave_awuser                                          (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                                              .awuser
		.hps_0_f2h_axi_slave_awvalid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                                              .awvalid
		.hps_0_f2h_axi_slave_awready                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                                              .awready
		.hps_0_f2h_axi_slave_wid                                             (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                                              .wid
		.hps_0_f2h_axi_slave_wdata                                           (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                                              .wdata
		.hps_0_f2h_axi_slave_wstrb                                           (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                                              .wstrb
		.hps_0_f2h_axi_slave_wlast                                           (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                                              .wlast
		.hps_0_f2h_axi_slave_wvalid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                                              .wvalid
		.hps_0_f2h_axi_slave_wready                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                                              .wready
		.hps_0_f2h_axi_slave_bid                                             (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                                              .bid
		.hps_0_f2h_axi_slave_bresp                                           (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                                              .bresp
		.hps_0_f2h_axi_slave_bvalid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                                              .bvalid
		.hps_0_f2h_axi_slave_bready                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                                              .bready
		.hps_0_f2h_axi_slave_arid                                            (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                                              .arid
		.hps_0_f2h_axi_slave_araddr                                          (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                                              .araddr
		.hps_0_f2h_axi_slave_arlen                                           (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                                              .arlen
		.hps_0_f2h_axi_slave_arsize                                          (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                                              .arsize
		.hps_0_f2h_axi_slave_arburst                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                                              .arburst
		.hps_0_f2h_axi_slave_arlock                                          (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                                              .arlock
		.hps_0_f2h_axi_slave_arcache                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                                              .arcache
		.hps_0_f2h_axi_slave_arprot                                          (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                                              .arprot
		.hps_0_f2h_axi_slave_aruser                                          (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                                              .aruser
		.hps_0_f2h_axi_slave_arvalid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                                              .arvalid
		.hps_0_f2h_axi_slave_arready                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                                              .arready
		.hps_0_f2h_axi_slave_rid                                             (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                                              .rid
		.hps_0_f2h_axi_slave_rdata                                           (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                                              .rdata
		.hps_0_f2h_axi_slave_rresp                                           (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                                              .rresp
		.hps_0_f2h_axi_slave_rlast                                           (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                                              .rlast
		.hps_0_f2h_axi_slave_rvalid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                                              .rvalid
		.hps_0_f2h_axi_slave_rready                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                       //                                                     clk_0_clk.clk
		.system_pll_outclk0_clk                                              (system_pll_outclk0_clk),                        //                                            system_pll_outclk0.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset    (rst_controller_005_reset_out_reset),            //    hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.hps_only_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                //               hps_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // hps_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_address                                      (hps_only_master_master_address),                //                                        hps_only_master_master.address
		.hps_only_master_master_waitrequest                                  (hps_only_master_master_waitrequest),            //                                                              .waitrequest
		.hps_only_master_master_byteenable                                   (hps_only_master_master_byteenable),             //                                                              .byteenable
		.hps_only_master_master_read                                         (hps_only_master_master_read),                   //                                                              .read
		.hps_only_master_master_readdata                                     (hps_only_master_master_readdata),               //                                                              .readdata
		.hps_only_master_master_readdatavalid                                (hps_only_master_master_readdatavalid),          //                                                              .readdatavalid
		.hps_only_master_master_write                                        (hps_only_master_master_write),                  //                                                              .write
		.hps_only_master_master_writedata                                    (hps_only_master_master_writedata)               //                                                              .writedata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.system_pll_outclk0_clk                                 (system_pll_outclk0_clk),                                    //                               system_pll_outclk0.clk
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.intr_capturer_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // intr_capturer_0_reset_sink_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                        (fpga_only_master_master_address),                           //                          fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                    (fpga_only_master_master_waitrequest),                       //                                                 .waitrequest
		.fpga_only_master_master_byteenable                     (fpga_only_master_master_byteenable),                        //                                                 .byteenable
		.fpga_only_master_master_read                           (fpga_only_master_master_read),                              //                                                 .read
		.fpga_only_master_master_readdata                       (fpga_only_master_master_readdata),                          //                                                 .readdata
		.fpga_only_master_master_readdatavalid                  (fpga_only_master_master_readdatavalid),                     //                                                 .readdatavalid
		.fpga_only_master_master_write                          (fpga_only_master_master_write),                             //                                                 .write
		.fpga_only_master_master_writedata                      (fpga_only_master_master_writedata),                         //                                                 .writedata
		.intr_capturer_0_avalon_slave_0_address                 (mm_interconnect_1_intr_capturer_0_avalon_slave_0_address),  //                   intr_capturer_0_avalon_slave_0.address
		.intr_capturer_0_avalon_slave_0_read                    (mm_interconnect_1_intr_capturer_0_avalon_slave_0_read),     //                                                 .read
		.intr_capturer_0_avalon_slave_0_readdata                (mm_interconnect_1_intr_capturer_0_avalon_slave_0_readdata), //                                                 .readdata
		.sysid_qsys_control_slave_address                       (mm_interconnect_1_sysid_qsys_control_slave_address),        //                         sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                      (mm_interconnect_1_sysid_qsys_control_slave_readdata)        //                                                 .readdata
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.system_pll_outclk0_clk                      (system_pll_outclk0_clk),                                        //                   system_pll_outclk0.clk
		.cpu_s0_reset_n_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                // cpu_s0_reset_n_reset_bridge_in_reset.reset
		.cpu_s0_data_master_address                  (cpu_s0_data_master_address),                                    //                   cpu_s0_data_master.address
		.cpu_s0_data_master_waitrequest              (cpu_s0_data_master_waitrequest),                                //                                     .waitrequest
		.cpu_s0_data_master_byteenable               (cpu_s0_data_master_byteenable),                                 //                                     .byteenable
		.cpu_s0_data_master_read                     (cpu_s0_data_master_read),                                       //                                     .read
		.cpu_s0_data_master_readdata                 (cpu_s0_data_master_readdata),                                   //                                     .readdata
		.cpu_s0_data_master_write                    (cpu_s0_data_master_write),                                      //                                     .write
		.cpu_s0_data_master_writedata                (cpu_s0_data_master_writedata),                                  //                                     .writedata
		.cpu_s0_data_master_debugaccess              (cpu_s0_data_master_debugaccess),                                //                                     .debugaccess
		.cpu_s0_instruction_master_address           (cpu_s0_instruction_master_address),                             //            cpu_s0_instruction_master.address
		.cpu_s0_instruction_master_waitrequest       (cpu_s0_instruction_master_waitrequest),                         //                                     .waitrequest
		.cpu_s0_instruction_master_burstcount        (cpu_s0_instruction_master_burstcount),                          //                                     .burstcount
		.cpu_s0_instruction_master_read              (cpu_s0_instruction_master_read),                                //                                     .read
		.cpu_s0_instruction_master_readdata          (cpu_s0_instruction_master_readdata),                            //                                     .readdata
		.cpu_s0_instruction_master_readdatavalid     (cpu_s0_instruction_master_readdatavalid),                       //                                     .readdatavalid
		.cpu_s0_jtag_debug_module_address            (mm_interconnect_2_cpu_s0_jtag_debug_module_address),            //             cpu_s0_jtag_debug_module.address
		.cpu_s0_jtag_debug_module_write              (mm_interconnect_2_cpu_s0_jtag_debug_module_write),              //                                     .write
		.cpu_s0_jtag_debug_module_read               (mm_interconnect_2_cpu_s0_jtag_debug_module_read),               //                                     .read
		.cpu_s0_jtag_debug_module_readdata           (mm_interconnect_2_cpu_s0_jtag_debug_module_readdata),           //                                     .readdata
		.cpu_s0_jtag_debug_module_writedata          (mm_interconnect_2_cpu_s0_jtag_debug_module_writedata),          //                                     .writedata
		.cpu_s0_jtag_debug_module_byteenable         (mm_interconnect_2_cpu_s0_jtag_debug_module_byteenable),         //                                     .byteenable
		.cpu_s0_jtag_debug_module_waitrequest        (mm_interconnect_2_cpu_s0_jtag_debug_module_waitrequest),        //                                     .waitrequest
		.cpu_s0_jtag_debug_module_debugaccess        (mm_interconnect_2_cpu_s0_jtag_debug_module_debugaccess),        //                                     .debugaccess
		.fifo_bridge_cpuM_cpus0_s0_address           (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_address),           //            fifo_bridge_cpuM_cpus0_s0.address
		.fifo_bridge_cpuM_cpus0_s0_write             (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_write),             //                                     .write
		.fifo_bridge_cpuM_cpus0_s0_read              (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_read),              //                                     .read
		.fifo_bridge_cpuM_cpus0_s0_readdata          (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_readdata),          //                                     .readdata
		.fifo_bridge_cpuM_cpus0_s0_writedata         (mm_interconnect_2_fifo_bridge_cpum_cpus0_s0_writedata),         //                                     .writedata
		.fifo_bridge_cpus0_cpus1_s0_address          (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_address),          //           fifo_bridge_cpus0_cpus1_s0.address
		.fifo_bridge_cpus0_cpus1_s0_write            (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_write),            //                                     .write
		.fifo_bridge_cpus0_cpus1_s0_read             (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_read),             //                                     .read
		.fifo_bridge_cpus0_cpus1_s0_readdata         (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_readdata),         //                                     .readdata
		.fifo_bridge_cpus0_cpus1_s0_writedata        (mm_interconnect_2_fifo_bridge_cpus0_cpus1_s0_writedata),        //                                     .writedata
		.s0_io_clockCrossing_bridge_s0_address       (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_address),       //        s0_io_clockCrossing_bridge_s0.address
		.s0_io_clockCrossing_bridge_s0_write         (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_write),         //                                     .write
		.s0_io_clockCrossing_bridge_s0_read          (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_read),          //                                     .read
		.s0_io_clockCrossing_bridge_s0_readdata      (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_readdata),      //                                     .readdata
		.s0_io_clockCrossing_bridge_s0_writedata     (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_writedata),     //                                     .writedata
		.s0_io_clockCrossing_bridge_s0_burstcount    (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_burstcount),    //                                     .burstcount
		.s0_io_clockCrossing_bridge_s0_byteenable    (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_byteenable),    //                                     .byteenable
		.s0_io_clockCrossing_bridge_s0_readdatavalid (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_readdatavalid), //                                     .readdatavalid
		.s0_io_clockCrossing_bridge_s0_waitrequest   (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_waitrequest),   //                                     .waitrequest
		.s0_io_clockCrossing_bridge_s0_debugaccess   (mm_interconnect_2_s0_io_clockcrossing_bridge_s0_debugaccess),   //                                     .debugaccess
		.sdram_clockCrossing_Bridge_s0_address       (mm_interconnect_2_sdram_clockcrossing_bridge_s0_address),       //        sdram_clockCrossing_Bridge_s0.address
		.sdram_clockCrossing_Bridge_s0_write         (mm_interconnect_2_sdram_clockcrossing_bridge_s0_write),         //                                     .write
		.sdram_clockCrossing_Bridge_s0_read          (mm_interconnect_2_sdram_clockcrossing_bridge_s0_read),          //                                     .read
		.sdram_clockCrossing_Bridge_s0_readdata      (mm_interconnect_2_sdram_clockcrossing_bridge_s0_readdata),      //                                     .readdata
		.sdram_clockCrossing_Bridge_s0_writedata     (mm_interconnect_2_sdram_clockcrossing_bridge_s0_writedata),     //                                     .writedata
		.sdram_clockCrossing_Bridge_s0_burstcount    (mm_interconnect_2_sdram_clockcrossing_bridge_s0_burstcount),    //                                     .burstcount
		.sdram_clockCrossing_Bridge_s0_byteenable    (mm_interconnect_2_sdram_clockcrossing_bridge_s0_byteenable),    //                                     .byteenable
		.sdram_clockCrossing_Bridge_s0_readdatavalid (mm_interconnect_2_sdram_clockcrossing_bridge_s0_readdatavalid), //                                     .readdatavalid
		.sdram_clockCrossing_Bridge_s0_waitrequest   (mm_interconnect_2_sdram_clockcrossing_bridge_s0_waitrequest),   //                                     .waitrequest
		.sdram_clockCrossing_Bridge_s0_debugaccess   (mm_interconnect_2_sdram_clockcrossing_bridge_s0_debugaccess)    //                                     .debugaccess
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                          //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                        //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                         //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                        //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                       //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                        //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                       //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                        //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                       //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                       //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                           //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                         //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                         //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                         //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                        //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                        //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                           //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                         //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                        //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                        //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                          //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                        //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                         //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                        //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                       //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                        //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                       //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                        //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                       //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                       //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                           //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                         //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                         //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                         //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                        //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                        //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                               //                                                     clk_0_clk.clk
		.system_pll_outclk0_clk                                              (system_pll_outclk0_clk),                                //                                            system_pll_outclk0.clk
		.fifo_bridge_cpuM_cpus0_clock_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                        //      fifo_bridge_cpuM_cpus0_clock_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                    // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.fifo_bridge_cpuM_cpus0_s1_address                                   (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_address),   //                                     fifo_bridge_cpuM_cpus0_s1.address
		.fifo_bridge_cpuM_cpus0_s1_write                                     (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_write),     //                                                              .write
		.fifo_bridge_cpuM_cpus0_s1_read                                      (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_read),      //                                                              .read
		.fifo_bridge_cpuM_cpus0_s1_readdata                                  (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_readdata),  //                                                              .readdata
		.fifo_bridge_cpuM_cpus0_s1_writedata                                 (mm_interconnect_3_fifo_bridge_cpum_cpus0_s1_writedata), //                                                              .writedata
		.fifo_bridge_cpuM_cpus1_s1_address                                   (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_address),   //                                     fifo_bridge_cpuM_cpus1_s1.address
		.fifo_bridge_cpuM_cpus1_s1_write                                     (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_write),     //                                                              .write
		.fifo_bridge_cpuM_cpus1_s1_read                                      (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_read),      //                                                              .read
		.fifo_bridge_cpuM_cpus1_s1_readdata                                  (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_readdata),  //                                                              .readdata
		.fifo_bridge_cpuM_cpus1_s1_writedata                                 (mm_interconnect_3_fifo_bridge_cpum_cpus1_s1_writedata)  //                                                              .writedata
	);

	soc_system_mm_interconnect_4 mm_interconnect_4 (
		.system_pll_outclk0_clk                      (system_pll_outclk0_clk),                                        //                   system_pll_outclk0.clk
		.cpu_s1_reset_n_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                // cpu_s1_reset_n_reset_bridge_in_reset.reset
		.cpu_s1_data_master_address                  (cpu_s1_data_master_address),                                    //                   cpu_s1_data_master.address
		.cpu_s1_data_master_waitrequest              (cpu_s1_data_master_waitrequest),                                //                                     .waitrequest
		.cpu_s1_data_master_byteenable               (cpu_s1_data_master_byteenable),                                 //                                     .byteenable
		.cpu_s1_data_master_read                     (cpu_s1_data_master_read),                                       //                                     .read
		.cpu_s1_data_master_readdata                 (cpu_s1_data_master_readdata),                                   //                                     .readdata
		.cpu_s1_data_master_write                    (cpu_s1_data_master_write),                                      //                                     .write
		.cpu_s1_data_master_writedata                (cpu_s1_data_master_writedata),                                  //                                     .writedata
		.cpu_s1_data_master_debugaccess              (cpu_s1_data_master_debugaccess),                                //                                     .debugaccess
		.cpu_s1_instruction_master_address           (cpu_s1_instruction_master_address),                             //            cpu_s1_instruction_master.address
		.cpu_s1_instruction_master_waitrequest       (cpu_s1_instruction_master_waitrequest),                         //                                     .waitrequest
		.cpu_s1_instruction_master_read              (cpu_s1_instruction_master_read),                                //                                     .read
		.cpu_s1_instruction_master_readdata          (cpu_s1_instruction_master_readdata),                            //                                     .readdata
		.cpu_s1_instruction_master_readdatavalid     (cpu_s1_instruction_master_readdatavalid),                       //                                     .readdatavalid
		.cpu_s1_jtag_debug_module_address            (mm_interconnect_4_cpu_s1_jtag_debug_module_address),            //             cpu_s1_jtag_debug_module.address
		.cpu_s1_jtag_debug_module_write              (mm_interconnect_4_cpu_s1_jtag_debug_module_write),              //                                     .write
		.cpu_s1_jtag_debug_module_read               (mm_interconnect_4_cpu_s1_jtag_debug_module_read),               //                                     .read
		.cpu_s1_jtag_debug_module_readdata           (mm_interconnect_4_cpu_s1_jtag_debug_module_readdata),           //                                     .readdata
		.cpu_s1_jtag_debug_module_writedata          (mm_interconnect_4_cpu_s1_jtag_debug_module_writedata),          //                                     .writedata
		.cpu_s1_jtag_debug_module_byteenable         (mm_interconnect_4_cpu_s1_jtag_debug_module_byteenable),         //                                     .byteenable
		.cpu_s1_jtag_debug_module_waitrequest        (mm_interconnect_4_cpu_s1_jtag_debug_module_waitrequest),        //                                     .waitrequest
		.cpu_s1_jtag_debug_module_debugaccess        (mm_interconnect_4_cpu_s1_jtag_debug_module_debugaccess),        //                                     .debugaccess
		.fifo_bridge_cpuM_cpus1_s0_address           (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_address),           //            fifo_bridge_cpuM_cpus1_s0.address
		.fifo_bridge_cpuM_cpus1_s0_write             (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_write),             //                                     .write
		.fifo_bridge_cpuM_cpus1_s0_read              (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_read),              //                                     .read
		.fifo_bridge_cpuM_cpus1_s0_readdata          (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_readdata),          //                                     .readdata
		.fifo_bridge_cpuM_cpus1_s0_writedata         (mm_interconnect_4_fifo_bridge_cpum_cpus1_s0_writedata),         //                                     .writedata
		.fifo_bridge_cpus0_cpus1_s1_address          (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_address),          //           fifo_bridge_cpus0_cpus1_s1.address
		.fifo_bridge_cpus0_cpus1_s1_write            (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_write),            //                                     .write
		.fifo_bridge_cpus0_cpus1_s1_read             (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_read),             //                                     .read
		.fifo_bridge_cpus0_cpus1_s1_readdata         (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_readdata),         //                                     .readdata
		.fifo_bridge_cpus0_cpus1_s1_writedata        (mm_interconnect_4_fifo_bridge_cpus0_cpus1_s1_writedata),        //                                     .writedata
		.onchip_sram_s1_address                      (mm_interconnect_4_onchip_sram_s1_address),                      //                       onchip_sram_s1.address
		.onchip_sram_s1_write                        (mm_interconnect_4_onchip_sram_s1_write),                        //                                     .write
		.onchip_sram_s1_readdata                     (mm_interconnect_4_onchip_sram_s1_readdata),                     //                                     .readdata
		.onchip_sram_s1_writedata                    (mm_interconnect_4_onchip_sram_s1_writedata),                    //                                     .writedata
		.onchip_sram_s1_byteenable                   (mm_interconnect_4_onchip_sram_s1_byteenable),                   //                                     .byteenable
		.onchip_sram_s1_chipselect                   (mm_interconnect_4_onchip_sram_s1_chipselect),                   //                                     .chipselect
		.onchip_sram_s1_clken                        (mm_interconnect_4_onchip_sram_s1_clken),                        //                                     .clken
		.s1_io_clockCrossing_bridge_s0_address       (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_address),       //        s1_io_clockCrossing_bridge_s0.address
		.s1_io_clockCrossing_bridge_s0_write         (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_write),         //                                     .write
		.s1_io_clockCrossing_bridge_s0_read          (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_read),          //                                     .read
		.s1_io_clockCrossing_bridge_s0_readdata      (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_readdata),      //                                     .readdata
		.s1_io_clockCrossing_bridge_s0_writedata     (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_writedata),     //                                     .writedata
		.s1_io_clockCrossing_bridge_s0_burstcount    (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_burstcount),    //                                     .burstcount
		.s1_io_clockCrossing_bridge_s0_byteenable    (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_byteenable),    //                                     .byteenable
		.s1_io_clockCrossing_bridge_s0_readdatavalid (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_readdatavalid), //                                     .readdatavalid
		.s1_io_clockCrossing_bridge_s0_waitrequest   (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_waitrequest),   //                                     .waitrequest
		.s1_io_clockCrossing_bridge_s0_debugaccess   (mm_interconnect_4_s1_io_clockcrossing_bridge_s0_debugaccess)    //                                     .debugaccess
	);

	soc_system_mm_interconnect_5 mm_interconnect_5 (
		.pwm_pll_outclk0_clk                                             (pwm_pll_outclk0_clk),                                              //                                           pwm_pll_outclk0.clk
		.system_pll_outclk1_clk                                          (system_pll_outclk1_clk),                                           //                                        system_pll_outclk1.clk
		.pwm_cpu_s0_1_clock_reset_reset_bridge_in_reset_reset            (rst_controller_004_reset_out_reset),                               //            pwm_cpu_s0_1_clock_reset_reset_bridge_in_reset.reset
		.s0_io_clockCrossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                               // s0_io_clockCrossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.s0_io_clockCrossing_bridge_m0_address                           (s0_io_clockcrossing_bridge_m0_address),                            //                             s0_io_clockCrossing_bridge_m0.address
		.s0_io_clockCrossing_bridge_m0_waitrequest                       (s0_io_clockcrossing_bridge_m0_waitrequest),                        //                                                          .waitrequest
		.s0_io_clockCrossing_bridge_m0_burstcount                        (s0_io_clockcrossing_bridge_m0_burstcount),                         //                                                          .burstcount
		.s0_io_clockCrossing_bridge_m0_byteenable                        (s0_io_clockcrossing_bridge_m0_byteenable),                         //                                                          .byteenable
		.s0_io_clockCrossing_bridge_m0_read                              (s0_io_clockcrossing_bridge_m0_read),                               //                                                          .read
		.s0_io_clockCrossing_bridge_m0_readdata                          (s0_io_clockcrossing_bridge_m0_readdata),                           //                                                          .readdata
		.s0_io_clockCrossing_bridge_m0_readdatavalid                     (s0_io_clockcrossing_bridge_m0_readdatavalid),                      //                                                          .readdatavalid
		.s0_io_clockCrossing_bridge_m0_write                             (s0_io_clockcrossing_bridge_m0_write),                              //                                                          .write
		.s0_io_clockCrossing_bridge_m0_writedata                         (s0_io_clockcrossing_bridge_m0_writedata),                          //                                                          .writedata
		.s0_io_clockCrossing_bridge_m0_debugaccess                       (s0_io_clockcrossing_bridge_m0_debugaccess),                        //                                                          .debugaccess
		.i2c_cpu_s0_mm_slave_address                                     (mm_interconnect_5_i2c_cpu_s0_mm_slave_address),                    //                                       i2c_cpu_s0_mm_slave.address
		.i2c_cpu_s0_mm_slave_write                                       (mm_interconnect_5_i2c_cpu_s0_mm_slave_write),                      //                                                          .write
		.i2c_cpu_s0_mm_slave_readdata                                    (mm_interconnect_5_i2c_cpu_s0_mm_slave_readdata),                   //                                                          .readdata
		.i2c_cpu_s0_mm_slave_writedata                                   (mm_interconnect_5_i2c_cpu_s0_mm_slave_writedata),                  //                                                          .writedata
		.i2c_cpu_s0_mm_slave_waitrequest                                 (~mm_interconnect_5_i2c_cpu_s0_mm_slave_waitrequest),               //                                                          .waitrequest
		.i2c_cpu_s0_mm_slave_chipselect                                  (mm_interconnect_5_i2c_cpu_s0_mm_slave_chipselect),                 //                                                          .chipselect
		.jtag_uart_cpu_s0_avalon_jtag_slave_address                      (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_address),     //                        jtag_uart_cpu_s0_avalon_jtag_slave.address
		.jtag_uart_cpu_s0_avalon_jtag_slave_write                        (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_write),       //                                                          .write
		.jtag_uart_cpu_s0_avalon_jtag_slave_read                         (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_read),        //                                                          .read
		.jtag_uart_cpu_s0_avalon_jtag_slave_readdata                     (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_readdata),    //                                                          .readdata
		.jtag_uart_cpu_s0_avalon_jtag_slave_writedata                    (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_writedata),   //                                                          .writedata
		.jtag_uart_cpu_s0_avalon_jtag_slave_waitrequest                  (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_waitrequest), //                                                          .waitrequest
		.jtag_uart_cpu_s0_avalon_jtag_slave_chipselect                   (mm_interconnect_5_jtag_uart_cpu_s0_avalon_jtag_slave_chipselect),  //                                                          .chipselect
		.pio_aliveTest_cpu_s0_s1_address                                 (mm_interconnect_5_pio_alivetest_cpu_s0_s1_address),                //                                   pio_aliveTest_cpu_s0_s1.address
		.pio_aliveTest_cpu_s0_s1_write                                   (mm_interconnect_5_pio_alivetest_cpu_s0_s1_write),                  //                                                          .write
		.pio_aliveTest_cpu_s0_s1_readdata                                (mm_interconnect_5_pio_alivetest_cpu_s0_s1_readdata),               //                                                          .readdata
		.pio_aliveTest_cpu_s0_s1_writedata                               (mm_interconnect_5_pio_alivetest_cpu_s0_s1_writedata),              //                                                          .writedata
		.pio_aliveTest_cpu_s0_s1_chipselect                              (mm_interconnect_5_pio_alivetest_cpu_s0_s1_chipselect),             //                                                          .chipselect
		.pwm_cpu_s0_1_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_1_s0_write),                          //                                           pwm_cpu_s0_1_s0.write
		.pwm_cpu_s0_1_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_1_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_2_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_2_s0_write),                          //                                           pwm_cpu_s0_2_s0.write
		.pwm_cpu_s0_2_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_2_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_3_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_3_s0_write),                          //                                           pwm_cpu_s0_3_s0.write
		.pwm_cpu_s0_3_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_3_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_4_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_4_s0_write),                          //                                           pwm_cpu_s0_4_s0.write
		.pwm_cpu_s0_4_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_4_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_5_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_5_s0_write),                          //                                           pwm_cpu_s0_5_s0.write
		.pwm_cpu_s0_5_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_5_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_6_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_6_s0_write),                          //                                           pwm_cpu_s0_6_s0.write
		.pwm_cpu_s0_6_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_6_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_7_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_7_s0_write),                          //                                           pwm_cpu_s0_7_s0.write
		.pwm_cpu_s0_7_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_7_s0_writedata),                      //                                                          .writedata
		.pwm_cpu_s0_8_s0_write                                           (mm_interconnect_5_pwm_cpu_s0_8_s0_write),                          //                                           pwm_cpu_s0_8_s0.write
		.pwm_cpu_s0_8_s0_writedata                                       (mm_interconnect_5_pwm_cpu_s0_8_s0_writedata),                      //                                                          .writedata
		.timer_cpu_s0_s1_address                                         (mm_interconnect_5_timer_cpu_s0_s1_address),                        //                                           timer_cpu_s0_s1.address
		.timer_cpu_s0_s1_write                                           (mm_interconnect_5_timer_cpu_s0_s1_write),                          //                                                          .write
		.timer_cpu_s0_s1_readdata                                        (mm_interconnect_5_timer_cpu_s0_s1_readdata),                       //                                                          .readdata
		.timer_cpu_s0_s1_writedata                                       (mm_interconnect_5_timer_cpu_s0_s1_writedata),                      //                                                          .writedata
		.timer_cpu_s0_s1_chipselect                                      (mm_interconnect_5_timer_cpu_s0_s1_chipselect)                      //                                                          .chipselect
	);

	soc_system_mm_interconnect_6 mm_interconnect_6 (
		.sdram_pll_outclk0_clk                                           (sdram_pll_outclk0_clk),                       //                                         sdram_pll_outclk0.clk
		.sdram_clockCrossing_Bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),          // sdram_clockCrossing_Bridge_m0_reset_reset_bridge_in_reset.reset
		.sdram_clockCrossing_Bridge_m0_address                           (sdram_clockcrossing_bridge_m0_address),       //                             sdram_clockCrossing_Bridge_m0.address
		.sdram_clockCrossing_Bridge_m0_waitrequest                       (sdram_clockcrossing_bridge_m0_waitrequest),   //                                                          .waitrequest
		.sdram_clockCrossing_Bridge_m0_burstcount                        (sdram_clockcrossing_bridge_m0_burstcount),    //                                                          .burstcount
		.sdram_clockCrossing_Bridge_m0_byteenable                        (sdram_clockcrossing_bridge_m0_byteenable),    //                                                          .byteenable
		.sdram_clockCrossing_Bridge_m0_read                              (sdram_clockcrossing_bridge_m0_read),          //                                                          .read
		.sdram_clockCrossing_Bridge_m0_readdata                          (sdram_clockcrossing_bridge_m0_readdata),      //                                                          .readdata
		.sdram_clockCrossing_Bridge_m0_readdatavalid                     (sdram_clockcrossing_bridge_m0_readdatavalid), //                                                          .readdatavalid
		.sdram_clockCrossing_Bridge_m0_write                             (sdram_clockcrossing_bridge_m0_write),         //                                                          .write
		.sdram_clockCrossing_Bridge_m0_writedata                         (sdram_clockcrossing_bridge_m0_writedata),     //                                                          .writedata
		.sdram_clockCrossing_Bridge_m0_debugaccess                       (sdram_clockcrossing_bridge_m0_debugaccess),   //                                                          .debugaccess
		.sdram_s1_address                                                (mm_interconnect_6_sdram_s1_address),          //                                                  sdram_s1.address
		.sdram_s1_write                                                  (mm_interconnect_6_sdram_s1_write),            //                                                          .write
		.sdram_s1_read                                                   (mm_interconnect_6_sdram_s1_read),             //                                                          .read
		.sdram_s1_readdata                                               (mm_interconnect_6_sdram_s1_readdata),         //                                                          .readdata
		.sdram_s1_writedata                                              (mm_interconnect_6_sdram_s1_writedata),        //                                                          .writedata
		.sdram_s1_byteenable                                             (mm_interconnect_6_sdram_s1_byteenable),       //                                                          .byteenable
		.sdram_s1_readdatavalid                                          (mm_interconnect_6_sdram_s1_readdatavalid),    //                                                          .readdatavalid
		.sdram_s1_waitrequest                                            (mm_interconnect_6_sdram_s1_waitrequest),      //                                                          .waitrequest
		.sdram_s1_chipselect                                             (mm_interconnect_6_sdram_s1_chipselect)        //                                                          .chipselect
	);

	soc_system_mm_interconnect_7 mm_interconnect_7 (
		.system_pll_outclk1_clk                                          (system_pll_outclk1_clk),                                           //                                        system_pll_outclk1.clk
		.s1_io_clockCrossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                               // s1_io_clockCrossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.s1_io_clockCrossing_bridge_m0_address                           (s1_io_clockcrossing_bridge_m0_address),                            //                             s1_io_clockCrossing_bridge_m0.address
		.s1_io_clockCrossing_bridge_m0_waitrequest                       (s1_io_clockcrossing_bridge_m0_waitrequest),                        //                                                          .waitrequest
		.s1_io_clockCrossing_bridge_m0_burstcount                        (s1_io_clockcrossing_bridge_m0_burstcount),                         //                                                          .burstcount
		.s1_io_clockCrossing_bridge_m0_byteenable                        (s1_io_clockcrossing_bridge_m0_byteenable),                         //                                                          .byteenable
		.s1_io_clockCrossing_bridge_m0_read                              (s1_io_clockcrossing_bridge_m0_read),                               //                                                          .read
		.s1_io_clockCrossing_bridge_m0_readdata                          (s1_io_clockcrossing_bridge_m0_readdata),                           //                                                          .readdata
		.s1_io_clockCrossing_bridge_m0_readdatavalid                     (s1_io_clockcrossing_bridge_m0_readdatavalid),                      //                                                          .readdatavalid
		.s1_io_clockCrossing_bridge_m0_write                             (s1_io_clockcrossing_bridge_m0_write),                              //                                                          .write
		.s1_io_clockCrossing_bridge_m0_writedata                         (s1_io_clockcrossing_bridge_m0_writedata),                          //                                                          .writedata
		.s1_io_clockCrossing_bridge_m0_debugaccess                       (s1_io_clockcrossing_bridge_m0_debugaccess),                        //                                                          .debugaccess
		.i2c_cpu_s1_mm_slave_address                                     (mm_interconnect_7_i2c_cpu_s1_mm_slave_address),                    //                                       i2c_cpu_s1_mm_slave.address
		.i2c_cpu_s1_mm_slave_write                                       (mm_interconnect_7_i2c_cpu_s1_mm_slave_write),                      //                                                          .write
		.i2c_cpu_s1_mm_slave_readdata                                    (mm_interconnect_7_i2c_cpu_s1_mm_slave_readdata),                   //                                                          .readdata
		.i2c_cpu_s1_mm_slave_writedata                                   (mm_interconnect_7_i2c_cpu_s1_mm_slave_writedata),                  //                                                          .writedata
		.i2c_cpu_s1_mm_slave_waitrequest                                 (~mm_interconnect_7_i2c_cpu_s1_mm_slave_waitrequest),               //                                                          .waitrequest
		.i2c_cpu_s1_mm_slave_chipselect                                  (mm_interconnect_7_i2c_cpu_s1_mm_slave_chipselect),                 //                                                          .chipselect
		.jtag_uart_cpu_s1_avalon_jtag_slave_address                      (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_address),     //                        jtag_uart_cpu_s1_avalon_jtag_slave.address
		.jtag_uart_cpu_s1_avalon_jtag_slave_write                        (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_write),       //                                                          .write
		.jtag_uart_cpu_s1_avalon_jtag_slave_read                         (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_read),        //                                                          .read
		.jtag_uart_cpu_s1_avalon_jtag_slave_readdata                     (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_readdata),    //                                                          .readdata
		.jtag_uart_cpu_s1_avalon_jtag_slave_writedata                    (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_writedata),   //                                                          .writedata
		.jtag_uart_cpu_s1_avalon_jtag_slave_waitrequest                  (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_waitrequest), //                                                          .waitrequest
		.jtag_uart_cpu_s1_avalon_jtag_slave_chipselect                   (mm_interconnect_7_jtag_uart_cpu_s1_avalon_jtag_slave_chipselect),  //                                                          .chipselect
		.pio_aliveTest_cpu_s1_s1_address                                 (mm_interconnect_7_pio_alivetest_cpu_s1_s1_address),                //                                   pio_aliveTest_cpu_s1_s1.address
		.pio_aliveTest_cpu_s1_s1_write                                   (mm_interconnect_7_pio_alivetest_cpu_s1_s1_write),                  //                                                          .write
		.pio_aliveTest_cpu_s1_s1_readdata                                (mm_interconnect_7_pio_alivetest_cpu_s1_s1_readdata),               //                                                          .readdata
		.pio_aliveTest_cpu_s1_s1_writedata                               (mm_interconnect_7_pio_alivetest_cpu_s1_s1_writedata),              //                                                          .writedata
		.pio_aliveTest_cpu_s1_s1_chipselect                              (mm_interconnect_7_pio_alivetest_cpu_s1_s1_chipselect),             //                                                          .chipselect
		.timer_cpu_s1_s1_address                                         (mm_interconnect_7_timer_cpu_s1_s1_address),                        //                                           timer_cpu_s1_s1.address
		.timer_cpu_s1_s1_write                                           (mm_interconnect_7_timer_cpu_s1_s1_write),                          //                                                          .write
		.timer_cpu_s1_s1_readdata                                        (mm_interconnect_7_timer_cpu_s1_s1_readdata),                       //                                                          .readdata
		.timer_cpu_s1_s1_writedata                                       (mm_interconnect_7_timer_cpu_s1_s1_writedata),                      //                                                          .writedata
		.timer_cpu_s1_s1_chipselect                                      (mm_interconnect_7_timer_cpu_s1_s1_chipselect)                      //                                                          .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_irq_mapper_002 irq_mapper_002 (
		.clk           (system_pll_outclk0_clk),                 //       clk.clk
		.reset         (rst_controller_reset_out_reset),         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver1_irq),               // receiver0.irq
		.receiver1_irq (irq_mapper_receiver0_irq),               // receiver1.irq
		.sender_irq    (intr_capturer_0_interrupt_receiver_irq)  //    sender.irq
	);

	soc_system_irq_mapper_003 irq_mapper_003 (
		.clk           (system_pll_outclk0_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),   // receiver1.irq
		.receiver2_irq (irq_mapper_003_receiver2_irq),   // receiver2.irq
		.receiver3_irq (irq_mapper_003_receiver3_irq),   // receiver3.irq
		.receiver4_irq (irq_mapper_003_receiver4_irq),   // receiver4.irq
		.sender_irq    (cpu_s0_d_irq_irq)                //    sender.irq
	);

	soc_system_irq_mapper_003 irq_mapper_004 (
		.clk           (system_pll_outclk0_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_004_receiver1_irq),   // receiver1.irq
		.receiver2_irq (irq_mapper_004_receiver2_irq),   // receiver2.irq
		.receiver3_irq (irq_mapper_004_receiver3_irq),   // receiver3.irq
		.receiver4_irq (irq_mapper_004_receiver4_irq),   // receiver4.irq
		.sender_irq    (cpu_s1_d_irq_irq)                //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (system_pll_outclk1_clk),             //       receiver_clk.clk
		.sender_clk     (system_pll_outclk0_clk),             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_003_receiver0_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (system_pll_outclk1_clk),             //       receiver_clk.clk
		.sender_clk     (system_pll_outclk0_clk),             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_003_receiver1_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (system_pll_outclk1_clk),             //       receiver_clk.clk
		.sender_clk     (system_pll_outclk0_clk),             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_003_receiver4_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (system_pll_outclk1_clk),             //       receiver_clk.clk
		.sender_clk     (system_pll_outclk0_clk),             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_004_receiver0_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (system_pll_outclk1_clk),             //       receiver_clk.clk
		.sender_clk     (system_pll_outclk0_clk),             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_004_receiver1_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (system_pll_outclk1_clk),             //       receiver_clk.clk
		.sender_clk     (system_pll_outclk0_clk),             //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_004_receiver4_irq)        //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (system_pll_outclk0_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (system_pll_outclk1_clk),             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pwm_pll_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
